module adresPortArbit(
  input         clock,
  input         reset,
  input         io_regEn,
  input         io_in_0_valid,
  input         io_in_1_valid,
  input         io_in_2_valid,
  input         io_in_3_valid,
  input         io_in_4_valid,
  input         io_in_5_valid,
  input         io_in_6_valid,
  input         io_in_7_valid,
  input         io_in_8_valid,
  input         io_in_9_valid,
  input         io_in_10_valid,
  input         io_in_11_valid,
  input         io_in_12_valid,
  input         io_in_13_valid,
  input         io_in_14_valid,
  input         io_in_15_valid,
  input         io_dmaEn,
  output [31:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  dmaNext; // @[outPortArbit.scala 98:24]
  wire  _T = ~dmaNext; // @[outPortArbit.scala 99:25]
  wire  _T_1 = io_dmaEn & _T; // @[outPortArbit.scala 99:22]
  wire  _T_3 = _T_1 | reset; // @[outPortArbit.scala 99:35]
  reg [3:0] indexReg; // @[Reg.scala 27:20]
  wire  _T_273 = 4'hf == indexReg; // @[Mux.scala 80:60]
  wire [3:0] _T_230 = io_in_13_valid ? 4'hd : 4'he; // @[Mux.scala 47:69]
  wire [3:0] _T_231 = io_in_12_valid ? 4'hc : _T_230; // @[Mux.scala 47:69]
  wire [3:0] _T_232 = io_in_11_valid ? 4'hb : _T_231; // @[Mux.scala 47:69]
  wire [3:0] _T_233 = io_in_10_valid ? 4'ha : _T_232; // @[Mux.scala 47:69]
  wire [3:0] _T_234 = io_in_9_valid ? 4'h9 : _T_233; // @[Mux.scala 47:69]
  wire [3:0] _T_235 = io_in_8_valid ? 4'h8 : _T_234; // @[Mux.scala 47:69]
  wire [3:0] _T_236 = io_in_7_valid ? 4'h7 : _T_235; // @[Mux.scala 47:69]
  wire [3:0] _T_237 = io_in_6_valid ? 4'h6 : _T_236; // @[Mux.scala 47:69]
  wire [3:0] _T_238 = io_in_5_valid ? 4'h5 : _T_237; // @[Mux.scala 47:69]
  wire [3:0] _T_239 = io_in_4_valid ? 4'h4 : _T_238; // @[Mux.scala 47:69]
  wire [3:0] _T_240 = io_in_3_valid ? 4'h3 : _T_239; // @[Mux.scala 47:69]
  wire [3:0] _T_241 = io_in_2_valid ? 4'h2 : _T_240; // @[Mux.scala 47:69]
  wire [3:0] _T_242 = io_in_1_valid ? 4'h1 : _T_241; // @[Mux.scala 47:69]
  wire [3:0] _T_243 = io_in_0_valid ? 4'h0 : _T_242; // @[Mux.scala 47:69]
  wire [3:0] _T_244 = io_in_15_valid ? 4'hf : _T_243; // @[Mux.scala 47:69]
  wire  _T_271 = 4'he == indexReg; // @[Mux.scala 80:60]
  wire [3:0] _T_215 = io_in_12_valid ? 4'hc : 4'hd; // @[Mux.scala 47:69]
  wire [3:0] _T_216 = io_in_11_valid ? 4'hb : _T_215; // @[Mux.scala 47:69]
  wire [3:0] _T_217 = io_in_10_valid ? 4'ha : _T_216; // @[Mux.scala 47:69]
  wire [3:0] _T_218 = io_in_9_valid ? 4'h9 : _T_217; // @[Mux.scala 47:69]
  wire [3:0] _T_219 = io_in_8_valid ? 4'h8 : _T_218; // @[Mux.scala 47:69]
  wire [3:0] _T_220 = io_in_7_valid ? 4'h7 : _T_219; // @[Mux.scala 47:69]
  wire [3:0] _T_221 = io_in_6_valid ? 4'h6 : _T_220; // @[Mux.scala 47:69]
  wire [3:0] _T_222 = io_in_5_valid ? 4'h5 : _T_221; // @[Mux.scala 47:69]
  wire [3:0] _T_223 = io_in_4_valid ? 4'h4 : _T_222; // @[Mux.scala 47:69]
  wire [3:0] _T_224 = io_in_3_valid ? 4'h3 : _T_223; // @[Mux.scala 47:69]
  wire [3:0] _T_225 = io_in_2_valid ? 4'h2 : _T_224; // @[Mux.scala 47:69]
  wire [3:0] _T_226 = io_in_1_valid ? 4'h1 : _T_225; // @[Mux.scala 47:69]
  wire [3:0] _T_227 = io_in_0_valid ? 4'h0 : _T_226; // @[Mux.scala 47:69]
  wire [3:0] _T_228 = io_in_15_valid ? 4'hf : _T_227; // @[Mux.scala 47:69]
  wire [3:0] _T_229 = io_in_14_valid ? 4'he : _T_228; // @[Mux.scala 47:69]
  wire  _T_269 = 4'hd == indexReg; // @[Mux.scala 80:60]
  wire [3:0] _T_200 = io_in_11_valid ? 4'hb : 4'hc; // @[Mux.scala 47:69]
  wire [3:0] _T_201 = io_in_10_valid ? 4'ha : _T_200; // @[Mux.scala 47:69]
  wire [3:0] _T_202 = io_in_9_valid ? 4'h9 : _T_201; // @[Mux.scala 47:69]
  wire [3:0] _T_203 = io_in_8_valid ? 4'h8 : _T_202; // @[Mux.scala 47:69]
  wire [3:0] _T_204 = io_in_7_valid ? 4'h7 : _T_203; // @[Mux.scala 47:69]
  wire [3:0] _T_205 = io_in_6_valid ? 4'h6 : _T_204; // @[Mux.scala 47:69]
  wire [3:0] _T_206 = io_in_5_valid ? 4'h5 : _T_205; // @[Mux.scala 47:69]
  wire [3:0] _T_207 = io_in_4_valid ? 4'h4 : _T_206; // @[Mux.scala 47:69]
  wire [3:0] _T_208 = io_in_3_valid ? 4'h3 : _T_207; // @[Mux.scala 47:69]
  wire [3:0] _T_209 = io_in_2_valid ? 4'h2 : _T_208; // @[Mux.scala 47:69]
  wire [3:0] _T_210 = io_in_1_valid ? 4'h1 : _T_209; // @[Mux.scala 47:69]
  wire [3:0] _T_211 = io_in_0_valid ? 4'h0 : _T_210; // @[Mux.scala 47:69]
  wire [3:0] _T_212 = io_in_15_valid ? 4'hf : _T_211; // @[Mux.scala 47:69]
  wire [3:0] _T_213 = io_in_14_valid ? 4'he : _T_212; // @[Mux.scala 47:69]
  wire [3:0] _T_214 = io_in_13_valid ? 4'hd : _T_213; // @[Mux.scala 47:69]
  wire  _T_267 = 4'hc == indexReg; // @[Mux.scala 80:60]
  wire [3:0] _T_185 = io_in_10_valid ? 4'ha : 4'hb; // @[Mux.scala 47:69]
  wire [3:0] _T_186 = io_in_9_valid ? 4'h9 : _T_185; // @[Mux.scala 47:69]
  wire [3:0] _T_187 = io_in_8_valid ? 4'h8 : _T_186; // @[Mux.scala 47:69]
  wire [3:0] _T_188 = io_in_7_valid ? 4'h7 : _T_187; // @[Mux.scala 47:69]
  wire [3:0] _T_189 = io_in_6_valid ? 4'h6 : _T_188; // @[Mux.scala 47:69]
  wire [3:0] _T_190 = io_in_5_valid ? 4'h5 : _T_189; // @[Mux.scala 47:69]
  wire [3:0] _T_191 = io_in_4_valid ? 4'h4 : _T_190; // @[Mux.scala 47:69]
  wire [3:0] _T_192 = io_in_3_valid ? 4'h3 : _T_191; // @[Mux.scala 47:69]
  wire [3:0] _T_193 = io_in_2_valid ? 4'h2 : _T_192; // @[Mux.scala 47:69]
  wire [3:0] _T_194 = io_in_1_valid ? 4'h1 : _T_193; // @[Mux.scala 47:69]
  wire [3:0] _T_195 = io_in_0_valid ? 4'h0 : _T_194; // @[Mux.scala 47:69]
  wire [3:0] _T_196 = io_in_15_valid ? 4'hf : _T_195; // @[Mux.scala 47:69]
  wire [3:0] _T_197 = io_in_14_valid ? 4'he : _T_196; // @[Mux.scala 47:69]
  wire [3:0] _T_198 = io_in_13_valid ? 4'hd : _T_197; // @[Mux.scala 47:69]
  wire [3:0] _T_199 = io_in_12_valid ? 4'hc : _T_198; // @[Mux.scala 47:69]
  wire  _T_265 = 4'hb == indexReg; // @[Mux.scala 80:60]
  wire [3:0] _T_170 = io_in_9_valid ? 4'h9 : 4'ha; // @[Mux.scala 47:69]
  wire [3:0] _T_171 = io_in_8_valid ? 4'h8 : _T_170; // @[Mux.scala 47:69]
  wire [3:0] _T_172 = io_in_7_valid ? 4'h7 : _T_171; // @[Mux.scala 47:69]
  wire [3:0] _T_173 = io_in_6_valid ? 4'h6 : _T_172; // @[Mux.scala 47:69]
  wire [3:0] _T_174 = io_in_5_valid ? 4'h5 : _T_173; // @[Mux.scala 47:69]
  wire [3:0] _T_175 = io_in_4_valid ? 4'h4 : _T_174; // @[Mux.scala 47:69]
  wire [3:0] _T_176 = io_in_3_valid ? 4'h3 : _T_175; // @[Mux.scala 47:69]
  wire [3:0] _T_177 = io_in_2_valid ? 4'h2 : _T_176; // @[Mux.scala 47:69]
  wire [3:0] _T_178 = io_in_1_valid ? 4'h1 : _T_177; // @[Mux.scala 47:69]
  wire [3:0] _T_179 = io_in_0_valid ? 4'h0 : _T_178; // @[Mux.scala 47:69]
  wire [3:0] _T_180 = io_in_15_valid ? 4'hf : _T_179; // @[Mux.scala 47:69]
  wire [3:0] _T_181 = io_in_14_valid ? 4'he : _T_180; // @[Mux.scala 47:69]
  wire [3:0] _T_182 = io_in_13_valid ? 4'hd : _T_181; // @[Mux.scala 47:69]
  wire [3:0] _T_183 = io_in_12_valid ? 4'hc : _T_182; // @[Mux.scala 47:69]
  wire [3:0] _T_184 = io_in_11_valid ? 4'hb : _T_183; // @[Mux.scala 47:69]
  wire  _T_263 = 4'ha == indexReg; // @[Mux.scala 80:60]
  wire [3:0] _T_155 = io_in_8_valid ? 4'h8 : 4'h9; // @[Mux.scala 47:69]
  wire [3:0] _T_156 = io_in_7_valid ? 4'h7 : _T_155; // @[Mux.scala 47:69]
  wire [3:0] _T_157 = io_in_6_valid ? 4'h6 : _T_156; // @[Mux.scala 47:69]
  wire [3:0] _T_158 = io_in_5_valid ? 4'h5 : _T_157; // @[Mux.scala 47:69]
  wire [3:0] _T_159 = io_in_4_valid ? 4'h4 : _T_158; // @[Mux.scala 47:69]
  wire [3:0] _T_160 = io_in_3_valid ? 4'h3 : _T_159; // @[Mux.scala 47:69]
  wire [3:0] _T_161 = io_in_2_valid ? 4'h2 : _T_160; // @[Mux.scala 47:69]
  wire [3:0] _T_162 = io_in_1_valid ? 4'h1 : _T_161; // @[Mux.scala 47:69]
  wire [3:0] _T_163 = io_in_0_valid ? 4'h0 : _T_162; // @[Mux.scala 47:69]
  wire [3:0] _T_164 = io_in_15_valid ? 4'hf : _T_163; // @[Mux.scala 47:69]
  wire [3:0] _T_165 = io_in_14_valid ? 4'he : _T_164; // @[Mux.scala 47:69]
  wire [3:0] _T_166 = io_in_13_valid ? 4'hd : _T_165; // @[Mux.scala 47:69]
  wire [3:0] _T_167 = io_in_12_valid ? 4'hc : _T_166; // @[Mux.scala 47:69]
  wire [3:0] _T_168 = io_in_11_valid ? 4'hb : _T_167; // @[Mux.scala 47:69]
  wire [3:0] _T_169 = io_in_10_valid ? 4'ha : _T_168; // @[Mux.scala 47:69]
  wire  _T_261 = 4'h9 == indexReg; // @[Mux.scala 80:60]
  wire [3:0] _T_140 = io_in_7_valid ? 4'h7 : 4'h8; // @[Mux.scala 47:69]
  wire [3:0] _T_141 = io_in_6_valid ? 4'h6 : _T_140; // @[Mux.scala 47:69]
  wire [3:0] _T_142 = io_in_5_valid ? 4'h5 : _T_141; // @[Mux.scala 47:69]
  wire [3:0] _T_143 = io_in_4_valid ? 4'h4 : _T_142; // @[Mux.scala 47:69]
  wire [3:0] _T_144 = io_in_3_valid ? 4'h3 : _T_143; // @[Mux.scala 47:69]
  wire [3:0] _T_145 = io_in_2_valid ? 4'h2 : _T_144; // @[Mux.scala 47:69]
  wire [3:0] _T_146 = io_in_1_valid ? 4'h1 : _T_145; // @[Mux.scala 47:69]
  wire [3:0] _T_147 = io_in_0_valid ? 4'h0 : _T_146; // @[Mux.scala 47:69]
  wire [3:0] _T_148 = io_in_15_valid ? 4'hf : _T_147; // @[Mux.scala 47:69]
  wire [3:0] _T_149 = io_in_14_valid ? 4'he : _T_148; // @[Mux.scala 47:69]
  wire [3:0] _T_150 = io_in_13_valid ? 4'hd : _T_149; // @[Mux.scala 47:69]
  wire [3:0] _T_151 = io_in_12_valid ? 4'hc : _T_150; // @[Mux.scala 47:69]
  wire [3:0] _T_152 = io_in_11_valid ? 4'hb : _T_151; // @[Mux.scala 47:69]
  wire [3:0] _T_153 = io_in_10_valid ? 4'ha : _T_152; // @[Mux.scala 47:69]
  wire [3:0] _T_154 = io_in_9_valid ? 4'h9 : _T_153; // @[Mux.scala 47:69]
  wire  _T_259 = 4'h8 == indexReg; // @[Mux.scala 80:60]
  wire [3:0] _T_125 = io_in_6_valid ? 4'h6 : 4'h7; // @[Mux.scala 47:69]
  wire [3:0] _T_126 = io_in_5_valid ? 4'h5 : _T_125; // @[Mux.scala 47:69]
  wire [3:0] _T_127 = io_in_4_valid ? 4'h4 : _T_126; // @[Mux.scala 47:69]
  wire [3:0] _T_128 = io_in_3_valid ? 4'h3 : _T_127; // @[Mux.scala 47:69]
  wire [3:0] _T_129 = io_in_2_valid ? 4'h2 : _T_128; // @[Mux.scala 47:69]
  wire [3:0] _T_130 = io_in_1_valid ? 4'h1 : _T_129; // @[Mux.scala 47:69]
  wire [3:0] _T_131 = io_in_0_valid ? 4'h0 : _T_130; // @[Mux.scala 47:69]
  wire [3:0] _T_132 = io_in_15_valid ? 4'hf : _T_131; // @[Mux.scala 47:69]
  wire [3:0] _T_133 = io_in_14_valid ? 4'he : _T_132; // @[Mux.scala 47:69]
  wire [3:0] _T_134 = io_in_13_valid ? 4'hd : _T_133; // @[Mux.scala 47:69]
  wire [3:0] _T_135 = io_in_12_valid ? 4'hc : _T_134; // @[Mux.scala 47:69]
  wire [3:0] _T_136 = io_in_11_valid ? 4'hb : _T_135; // @[Mux.scala 47:69]
  wire [3:0] _T_137 = io_in_10_valid ? 4'ha : _T_136; // @[Mux.scala 47:69]
  wire [3:0] _T_138 = io_in_9_valid ? 4'h9 : _T_137; // @[Mux.scala 47:69]
  wire [3:0] _T_139 = io_in_8_valid ? 4'h8 : _T_138; // @[Mux.scala 47:69]
  wire  _T_257 = 4'h7 == indexReg; // @[Mux.scala 80:60]
  wire [3:0] _T_110 = io_in_5_valid ? 4'h5 : 4'h6; // @[Mux.scala 47:69]
  wire [3:0] _T_111 = io_in_4_valid ? 4'h4 : _T_110; // @[Mux.scala 47:69]
  wire [3:0] _T_112 = io_in_3_valid ? 4'h3 : _T_111; // @[Mux.scala 47:69]
  wire [3:0] _T_113 = io_in_2_valid ? 4'h2 : _T_112; // @[Mux.scala 47:69]
  wire [3:0] _T_114 = io_in_1_valid ? 4'h1 : _T_113; // @[Mux.scala 47:69]
  wire [3:0] _T_115 = io_in_0_valid ? 4'h0 : _T_114; // @[Mux.scala 47:69]
  wire [3:0] _T_116 = io_in_15_valid ? 4'hf : _T_115; // @[Mux.scala 47:69]
  wire [3:0] _T_117 = io_in_14_valid ? 4'he : _T_116; // @[Mux.scala 47:69]
  wire [3:0] _T_118 = io_in_13_valid ? 4'hd : _T_117; // @[Mux.scala 47:69]
  wire [3:0] _T_119 = io_in_12_valid ? 4'hc : _T_118; // @[Mux.scala 47:69]
  wire [3:0] _T_120 = io_in_11_valid ? 4'hb : _T_119; // @[Mux.scala 47:69]
  wire [3:0] _T_121 = io_in_10_valid ? 4'ha : _T_120; // @[Mux.scala 47:69]
  wire [3:0] _T_122 = io_in_9_valid ? 4'h9 : _T_121; // @[Mux.scala 47:69]
  wire [3:0] _T_123 = io_in_8_valid ? 4'h8 : _T_122; // @[Mux.scala 47:69]
  wire [3:0] _T_124 = io_in_7_valid ? 4'h7 : _T_123; // @[Mux.scala 47:69]
  wire  _T_255 = 4'h6 == indexReg; // @[Mux.scala 80:60]
  wire [3:0] _T_95 = io_in_4_valid ? 4'h4 : 4'h5; // @[Mux.scala 47:69]
  wire [3:0] _T_96 = io_in_3_valid ? 4'h3 : _T_95; // @[Mux.scala 47:69]
  wire [3:0] _T_97 = io_in_2_valid ? 4'h2 : _T_96; // @[Mux.scala 47:69]
  wire [3:0] _T_98 = io_in_1_valid ? 4'h1 : _T_97; // @[Mux.scala 47:69]
  wire [3:0] _T_99 = io_in_0_valid ? 4'h0 : _T_98; // @[Mux.scala 47:69]
  wire [3:0] _T_100 = io_in_15_valid ? 4'hf : _T_99; // @[Mux.scala 47:69]
  wire [3:0] _T_101 = io_in_14_valid ? 4'he : _T_100; // @[Mux.scala 47:69]
  wire [3:0] _T_102 = io_in_13_valid ? 4'hd : _T_101; // @[Mux.scala 47:69]
  wire [3:0] _T_103 = io_in_12_valid ? 4'hc : _T_102; // @[Mux.scala 47:69]
  wire [3:0] _T_104 = io_in_11_valid ? 4'hb : _T_103; // @[Mux.scala 47:69]
  wire [3:0] _T_105 = io_in_10_valid ? 4'ha : _T_104; // @[Mux.scala 47:69]
  wire [3:0] _T_106 = io_in_9_valid ? 4'h9 : _T_105; // @[Mux.scala 47:69]
  wire [3:0] _T_107 = io_in_8_valid ? 4'h8 : _T_106; // @[Mux.scala 47:69]
  wire [3:0] _T_108 = io_in_7_valid ? 4'h7 : _T_107; // @[Mux.scala 47:69]
  wire [3:0] _T_109 = io_in_6_valid ? 4'h6 : _T_108; // @[Mux.scala 47:69]
  wire  _T_253 = 4'h5 == indexReg; // @[Mux.scala 80:60]
  wire [3:0] _T_80 = io_in_3_valid ? 4'h3 : 4'h4; // @[Mux.scala 47:69]
  wire [3:0] _T_81 = io_in_2_valid ? 4'h2 : _T_80; // @[Mux.scala 47:69]
  wire [3:0] _T_82 = io_in_1_valid ? 4'h1 : _T_81; // @[Mux.scala 47:69]
  wire [3:0] _T_83 = io_in_0_valid ? 4'h0 : _T_82; // @[Mux.scala 47:69]
  wire [3:0] _T_84 = io_in_15_valid ? 4'hf : _T_83; // @[Mux.scala 47:69]
  wire [3:0] _T_85 = io_in_14_valid ? 4'he : _T_84; // @[Mux.scala 47:69]
  wire [3:0] _T_86 = io_in_13_valid ? 4'hd : _T_85; // @[Mux.scala 47:69]
  wire [3:0] _T_87 = io_in_12_valid ? 4'hc : _T_86; // @[Mux.scala 47:69]
  wire [3:0] _T_88 = io_in_11_valid ? 4'hb : _T_87; // @[Mux.scala 47:69]
  wire [3:0] _T_89 = io_in_10_valid ? 4'ha : _T_88; // @[Mux.scala 47:69]
  wire [3:0] _T_90 = io_in_9_valid ? 4'h9 : _T_89; // @[Mux.scala 47:69]
  wire [3:0] _T_91 = io_in_8_valid ? 4'h8 : _T_90; // @[Mux.scala 47:69]
  wire [3:0] _T_92 = io_in_7_valid ? 4'h7 : _T_91; // @[Mux.scala 47:69]
  wire [3:0] _T_93 = io_in_6_valid ? 4'h6 : _T_92; // @[Mux.scala 47:69]
  wire [3:0] _T_94 = io_in_5_valid ? 4'h5 : _T_93; // @[Mux.scala 47:69]
  wire  _T_251 = 4'h4 == indexReg; // @[Mux.scala 80:60]
  wire [3:0] _T_65 = io_in_2_valid ? 4'h2 : 4'h3; // @[Mux.scala 47:69]
  wire [3:0] _T_66 = io_in_1_valid ? 4'h1 : _T_65; // @[Mux.scala 47:69]
  wire [3:0] _T_67 = io_in_0_valid ? 4'h0 : _T_66; // @[Mux.scala 47:69]
  wire [3:0] _T_68 = io_in_15_valid ? 4'hf : _T_67; // @[Mux.scala 47:69]
  wire [3:0] _T_69 = io_in_14_valid ? 4'he : _T_68; // @[Mux.scala 47:69]
  wire [3:0] _T_70 = io_in_13_valid ? 4'hd : _T_69; // @[Mux.scala 47:69]
  wire [3:0] _T_71 = io_in_12_valid ? 4'hc : _T_70; // @[Mux.scala 47:69]
  wire [3:0] _T_72 = io_in_11_valid ? 4'hb : _T_71; // @[Mux.scala 47:69]
  wire [3:0] _T_73 = io_in_10_valid ? 4'ha : _T_72; // @[Mux.scala 47:69]
  wire [3:0] _T_74 = io_in_9_valid ? 4'h9 : _T_73; // @[Mux.scala 47:69]
  wire [3:0] _T_75 = io_in_8_valid ? 4'h8 : _T_74; // @[Mux.scala 47:69]
  wire [3:0] _T_76 = io_in_7_valid ? 4'h7 : _T_75; // @[Mux.scala 47:69]
  wire [3:0] _T_77 = io_in_6_valid ? 4'h6 : _T_76; // @[Mux.scala 47:69]
  wire [3:0] _T_78 = io_in_5_valid ? 4'h5 : _T_77; // @[Mux.scala 47:69]
  wire [3:0] _T_79 = io_in_4_valid ? 4'h4 : _T_78; // @[Mux.scala 47:69]
  wire  _T_249 = 4'h3 == indexReg; // @[Mux.scala 80:60]
  wire [3:0] _T_50 = io_in_1_valid ? 4'h1 : 4'h2; // @[Mux.scala 47:69]
  wire [3:0] _T_51 = io_in_0_valid ? 4'h0 : _T_50; // @[Mux.scala 47:69]
  wire [3:0] _T_52 = io_in_15_valid ? 4'hf : _T_51; // @[Mux.scala 47:69]
  wire [3:0] _T_53 = io_in_14_valid ? 4'he : _T_52; // @[Mux.scala 47:69]
  wire [3:0] _T_54 = io_in_13_valid ? 4'hd : _T_53; // @[Mux.scala 47:69]
  wire [3:0] _T_55 = io_in_12_valid ? 4'hc : _T_54; // @[Mux.scala 47:69]
  wire [3:0] _T_56 = io_in_11_valid ? 4'hb : _T_55; // @[Mux.scala 47:69]
  wire [3:0] _T_57 = io_in_10_valid ? 4'ha : _T_56; // @[Mux.scala 47:69]
  wire [3:0] _T_58 = io_in_9_valid ? 4'h9 : _T_57; // @[Mux.scala 47:69]
  wire [3:0] _T_59 = io_in_8_valid ? 4'h8 : _T_58; // @[Mux.scala 47:69]
  wire [3:0] _T_60 = io_in_7_valid ? 4'h7 : _T_59; // @[Mux.scala 47:69]
  wire [3:0] _T_61 = io_in_6_valid ? 4'h6 : _T_60; // @[Mux.scala 47:69]
  wire [3:0] _T_62 = io_in_5_valid ? 4'h5 : _T_61; // @[Mux.scala 47:69]
  wire [3:0] _T_63 = io_in_4_valid ? 4'h4 : _T_62; // @[Mux.scala 47:69]
  wire [3:0] _T_64 = io_in_3_valid ? 4'h3 : _T_63; // @[Mux.scala 47:69]
  wire  _T_247 = 4'h2 == indexReg; // @[Mux.scala 80:60]
  wire [3:0] _T_35 = io_in_0_valid ? 4'h0 : 4'h1; // @[Mux.scala 47:69]
  wire [3:0] _T_36 = io_in_15_valid ? 4'hf : _T_35; // @[Mux.scala 47:69]
  wire [3:0] _T_37 = io_in_14_valid ? 4'he : _T_36; // @[Mux.scala 47:69]
  wire [3:0] _T_38 = io_in_13_valid ? 4'hd : _T_37; // @[Mux.scala 47:69]
  wire [3:0] _T_39 = io_in_12_valid ? 4'hc : _T_38; // @[Mux.scala 47:69]
  wire [3:0] _T_40 = io_in_11_valid ? 4'hb : _T_39; // @[Mux.scala 47:69]
  wire [3:0] _T_41 = io_in_10_valid ? 4'ha : _T_40; // @[Mux.scala 47:69]
  wire [3:0] _T_42 = io_in_9_valid ? 4'h9 : _T_41; // @[Mux.scala 47:69]
  wire [3:0] _T_43 = io_in_8_valid ? 4'h8 : _T_42; // @[Mux.scala 47:69]
  wire [3:0] _T_44 = io_in_7_valid ? 4'h7 : _T_43; // @[Mux.scala 47:69]
  wire [3:0] _T_45 = io_in_6_valid ? 4'h6 : _T_44; // @[Mux.scala 47:69]
  wire [3:0] _T_46 = io_in_5_valid ? 4'h5 : _T_45; // @[Mux.scala 47:69]
  wire [3:0] _T_47 = io_in_4_valid ? 4'h4 : _T_46; // @[Mux.scala 47:69]
  wire [3:0] _T_48 = io_in_3_valid ? 4'h3 : _T_47; // @[Mux.scala 47:69]
  wire [3:0] _T_49 = io_in_2_valid ? 4'h2 : _T_48; // @[Mux.scala 47:69]
  wire  _T_245 = 4'h1 == indexReg; // @[Mux.scala 80:60]
  wire [3:0] _T_20 = io_in_15_valid ? 4'hf : 4'h0; // @[Mux.scala 47:69]
  wire [3:0] _T_21 = io_in_14_valid ? 4'he : _T_20; // @[Mux.scala 47:69]
  wire [3:0] _T_22 = io_in_13_valid ? 4'hd : _T_21; // @[Mux.scala 47:69]
  wire [3:0] _T_23 = io_in_12_valid ? 4'hc : _T_22; // @[Mux.scala 47:69]
  wire [3:0] _T_24 = io_in_11_valid ? 4'hb : _T_23; // @[Mux.scala 47:69]
  wire [3:0] _T_25 = io_in_10_valid ? 4'ha : _T_24; // @[Mux.scala 47:69]
  wire [3:0] _T_26 = io_in_9_valid ? 4'h9 : _T_25; // @[Mux.scala 47:69]
  wire [3:0] _T_27 = io_in_8_valid ? 4'h8 : _T_26; // @[Mux.scala 47:69]
  wire [3:0] _T_28 = io_in_7_valid ? 4'h7 : _T_27; // @[Mux.scala 47:69]
  wire [3:0] _T_29 = io_in_6_valid ? 4'h6 : _T_28; // @[Mux.scala 47:69]
  wire [3:0] _T_30 = io_in_5_valid ? 4'h5 : _T_29; // @[Mux.scala 47:69]
  wire [3:0] _T_31 = io_in_4_valid ? 4'h4 : _T_30; // @[Mux.scala 47:69]
  wire [3:0] _T_32 = io_in_3_valid ? 4'h3 : _T_31; // @[Mux.scala 47:69]
  wire [3:0] _T_33 = io_in_2_valid ? 4'h2 : _T_32; // @[Mux.scala 47:69]
  wire [3:0] _T_34 = io_in_1_valid ? 4'h1 : _T_33; // @[Mux.scala 47:69]
  wire [3:0] _T_5 = io_in_14_valid ? 4'he : 4'hf; // @[Mux.scala 47:69]
  wire [3:0] _T_6 = io_in_13_valid ? 4'hd : _T_5; // @[Mux.scala 47:69]
  wire [3:0] _T_7 = io_in_12_valid ? 4'hc : _T_6; // @[Mux.scala 47:69]
  wire [3:0] _T_8 = io_in_11_valid ? 4'hb : _T_7; // @[Mux.scala 47:69]
  wire [3:0] _T_9 = io_in_10_valid ? 4'ha : _T_8; // @[Mux.scala 47:69]
  wire [3:0] _T_10 = io_in_9_valid ? 4'h9 : _T_9; // @[Mux.scala 47:69]
  wire [3:0] _T_11 = io_in_8_valid ? 4'h8 : _T_10; // @[Mux.scala 47:69]
  wire [3:0] _T_12 = io_in_7_valid ? 4'h7 : _T_11; // @[Mux.scala 47:69]
  wire [3:0] _T_13 = io_in_6_valid ? 4'h6 : _T_12; // @[Mux.scala 47:69]
  wire [3:0] _T_14 = io_in_5_valid ? 4'h5 : _T_13; // @[Mux.scala 47:69]
  wire [3:0] _T_15 = io_in_4_valid ? 4'h4 : _T_14; // @[Mux.scala 47:69]
  wire [3:0] _T_16 = io_in_3_valid ? 4'h3 : _T_15; // @[Mux.scala 47:69]
  wire [3:0] _T_17 = io_in_2_valid ? 4'h2 : _T_16; // @[Mux.scala 47:69]
  wire [3:0] _T_18 = io_in_1_valid ? 4'h1 : _T_17; // @[Mux.scala 47:69]
  wire [3:0] _T_19 = io_in_0_valid ? 4'h0 : _T_18; // @[Mux.scala 47:69]
  wire [3:0] _T_246 = _T_245 ? _T_34 : _T_19; // @[Mux.scala 80:57]
  wire [3:0] _T_248 = _T_247 ? _T_49 : _T_246; // @[Mux.scala 80:57]
  wire [3:0] _T_250 = _T_249 ? _T_64 : _T_248; // @[Mux.scala 80:57]
  wire [3:0] _T_252 = _T_251 ? _T_79 : _T_250; // @[Mux.scala 80:57]
  wire [3:0] _T_254 = _T_253 ? _T_94 : _T_252; // @[Mux.scala 80:57]
  wire [3:0] _T_256 = _T_255 ? _T_109 : _T_254; // @[Mux.scala 80:57]
  wire [3:0] _T_258 = _T_257 ? _T_124 : _T_256; // @[Mux.scala 80:57]
  wire [3:0] _T_260 = _T_259 ? _T_139 : _T_258; // @[Mux.scala 80:57]
  wire [3:0] _T_262 = _T_261 ? _T_154 : _T_260; // @[Mux.scala 80:57]
  wire [3:0] _T_264 = _T_263 ? _T_169 : _T_262; // @[Mux.scala 80:57]
  wire [3:0] _T_266 = _T_265 ? _T_184 : _T_264; // @[Mux.scala 80:57]
  wire [3:0] _T_268 = _T_267 ? _T_199 : _T_266; // @[Mux.scala 80:57]
  wire [3:0] _T_270 = _T_269 ? _T_214 : _T_268; // @[Mux.scala 80:57]
  wire [3:0] _T_272 = _T_271 ? _T_229 : _T_270; // @[Mux.scala 80:57]
  wire [3:0] selOut = _T_273 ? _T_244 : _T_272; // @[Mux.scala 80:57]
  wire [3:0] _T_275 = selOut + 4'h1; // @[outPortArbit.scala 117:27]
  wire [4:0] _GEN_2 = {{1'd0}, _T_275}; // @[outPortArbit.scala 117:34]
  wire  _T_276 = _GEN_2 == 5'h10; // @[outPortArbit.scala 117:34]
  wire  _T_280 = 4'h1 == selOut; // @[Mux.scala 80:60]
  wire  _T_282 = 4'h2 == selOut; // @[Mux.scala 80:60]
  wire  _T_284 = 4'h3 == selOut; // @[Mux.scala 80:60]
  wire  _T_286 = 4'h4 == selOut; // @[Mux.scala 80:60]
  wire  _T_288 = 4'h5 == selOut; // @[Mux.scala 80:60]
  wire  _T_290 = 4'h6 == selOut; // @[Mux.scala 80:60]
  wire  _T_292 = 4'h7 == selOut; // @[Mux.scala 80:60]
  wire  _T_294 = 4'h8 == selOut; // @[Mux.scala 80:60]
  wire  _T_296 = 4'h9 == selOut; // @[Mux.scala 80:60]
  wire  _T_298 = 4'ha == selOut; // @[Mux.scala 80:60]
  wire  _T_300 = 4'hb == selOut; // @[Mux.scala 80:60]
  wire  _T_302 = 4'hc == selOut; // @[Mux.scala 80:60]
  wire  _T_304 = 4'hd == selOut; // @[Mux.scala 80:60]
  wire  _T_306 = 4'he == selOut; // @[Mux.scala 80:60]
  wire  _T_308 = 4'hf == selOut; // @[Mux.scala 80:60]
  reg [31:0] _T_310; // @[Reg.scala 27:20]
  assign io_out = _T_310; // @[outPortArbit.scala 120:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dmaNext = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  indexReg = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  _T_310 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    dmaNext <= io_dmaEn;
    if (_T_3) begin
      indexReg <= 4'h0;
    end else if (io_regEn) begin
      if (_T_276) begin
        indexReg <= 4'h0;
      end else begin
        indexReg <= _T_275;
      end
    end
    if (reset) begin
      _T_310 <= 32'h0;
    end else if (io_regEn) begin
      if (_T_308) begin
        _T_310 <= 32'h201007c;
      end else if (_T_306) begin
        _T_310 <= 32'h2010078;
      end else if (_T_304) begin
        _T_310 <= 32'h2010074;
      end else if (_T_302) begin
        _T_310 <= 32'h2010070;
      end else if (_T_300) begin
        _T_310 <= 32'h201006c;
      end else if (_T_298) begin
        _T_310 <= 32'h2010068;
      end else if (_T_296) begin
        _T_310 <= 32'h2010064;
      end else if (_T_294) begin
        _T_310 <= 32'h2010060;
      end else if (_T_292) begin
        _T_310 <= 32'h201005c;
      end else if (_T_290) begin
        _T_310 <= 32'h2010058;
      end else if (_T_288) begin
        _T_310 <= 32'h2010054;
      end else if (_T_286) begin
        _T_310 <= 32'h2010050;
      end else if (_T_284) begin
        _T_310 <= 32'h201004c;
      end else if (_T_282) begin
        _T_310 <= 32'h2010048;
      end else if (_T_280) begin
        _T_310 <= 32'h2010044;
      end else begin
        _T_310 <= 32'h2010040;
      end
    end
  end
endmodule
module DMACtrl(
  input          clock,
  input          reset,
  input          io_dataIn_awready,
  output         io_dataIn_awvalid,
  output [31:0]  io_dataIn_awaddr,
  output [7:0]   io_dataIn_awlen,
  input          io_dataIn_wready,
  output         io_dataIn_wvalid,
  output [63:0]  io_dataIn_wdata,
  output         io_dataIn_wlast,
  output         io_dataIn_bready,
  input          io_dataIn_bvalid,
  input          io_dataIn_arready,
  output         io_dataIn_arvalid,
  output [31:0]  io_dataIn_araddr,
  output [7:0]   io_dataIn_arlen,
  output         io_dataIn_rready,
  input          io_dataIn_rvalid,
  input  [63:0]  io_dataIn_rdata,
  input          io_dataIn_rlast,
  output         io_dataOutMMIO_valid,
  input          io_dataOutMMIO_ready,
  input  [63:0]  io_dataOutMMIO_data_read,
  output [63:0]  io_dataOutMMIO_data_write,
  output         io_dataOutMMIO_wen,
  output [31:0]  io_dataOutMMIO_addr,
  input          dmaEn_0,
  input          dmaEnWR_0,
  input          block3_0,
  input  [191:0] dmaCtrl_0,
  input          block2_0,
  output         blockDMA_0,
  output         DMABuzy_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  portArbitInst_clock; // @[DMACtrlWRMask.scala 56:29]
  wire  portArbitInst_reset; // @[DMACtrlWRMask.scala 56:29]
  wire  portArbitInst_io_regEn; // @[DMACtrlWRMask.scala 56:29]
  wire  portArbitInst_io_in_0_valid; // @[DMACtrlWRMask.scala 56:29]
  wire  portArbitInst_io_in_1_valid; // @[DMACtrlWRMask.scala 56:29]
  wire  portArbitInst_io_in_2_valid; // @[DMACtrlWRMask.scala 56:29]
  wire  portArbitInst_io_in_3_valid; // @[DMACtrlWRMask.scala 56:29]
  wire  portArbitInst_io_in_4_valid; // @[DMACtrlWRMask.scala 56:29]
  wire  portArbitInst_io_in_5_valid; // @[DMACtrlWRMask.scala 56:29]
  wire  portArbitInst_io_in_6_valid; // @[DMACtrlWRMask.scala 56:29]
  wire  portArbitInst_io_in_7_valid; // @[DMACtrlWRMask.scala 56:29]
  wire  portArbitInst_io_in_8_valid; // @[DMACtrlWRMask.scala 56:29]
  wire  portArbitInst_io_in_9_valid; // @[DMACtrlWRMask.scala 56:29]
  wire  portArbitInst_io_in_10_valid; // @[DMACtrlWRMask.scala 56:29]
  wire  portArbitInst_io_in_11_valid; // @[DMACtrlWRMask.scala 56:29]
  wire  portArbitInst_io_in_12_valid; // @[DMACtrlWRMask.scala 56:29]
  wire  portArbitInst_io_in_13_valid; // @[DMACtrlWRMask.scala 56:29]
  wire  portArbitInst_io_in_14_valid; // @[DMACtrlWRMask.scala 56:29]
  wire  portArbitInst_io_in_15_valid; // @[DMACtrlWRMask.scala 56:29]
  wire  portArbitInst_io_dmaEn; // @[DMACtrlWRMask.scala 56:29]
  wire [31:0] portArbitInst_io_out; // @[DMACtrlWRMask.scala 56:29]
  wire  block = block2_0 | block3_0; // @[DMACtrlWRMask.scala 37:22]
  wire [31:0] dmaAXIAddrR = dmaCtrl_0[31:0]; // @[DMACtrlWRMask.scala 41:28]
  wire [31:0] dmaCGRAOutMask = dmaCtrl_0[127:96]; // @[DMACtrlWRMask.scala 44:31]
  wire [31:0] dmaLenR = dmaCtrl_0[159:128]; // @[DMACtrlWRMask.scala 45:24]
  wire [31:0] dmaLenW = dmaCtrl_0[191:160]; // @[DMACtrlWRMask.scala 46:24]
  wire [63:0] dmaAXIAddr = dmaCtrl_0[63:0]; // @[DMACtrlWRMask.scala 49:27]
  wire [63:0] dmaDstAddr = dmaCtrl_0[127:64]; // @[DMACtrlWRMask.scala 50:27]
  wire [63:0] dmaLen = dmaCtrl_0[191:128]; // @[DMACtrlWRMask.scala 51:23]
  wire  isCfg = dmaDstAddr == 64'h2010080; // @[DMACtrlWRMask.scala 52:26]
  reg  changeState; // @[DMACtrlWRMask.scala 75:28]
  reg [1:0] rState; // @[DMACtrlWRMask.scala 80:23]
  wire  _T_64 = dmaEn_0 | dmaEnWR_0; // @[DMACtrlWRMask.scala 81:31]
  reg  dmaNext; // @[DMACtrlWRMask.scala 81:24]
  wire  _T_66 = ~dmaNext; // @[DMACtrlWRMask.scala 82:42]
  wire  _T_67 = _T_64 & _T_66; // @[DMACtrlWRMask.scala 82:39]
  wire  _T_68 = ~changeState; // @[DMACtrlWRMask.scala 82:54]
  wire  _T_69 = _T_67 & _T_68; // @[DMACtrlWRMask.scala 82:51]
  wire  _T_71 = io_dataIn_arready & _T_68; // @[DMACtrlWRMask.scala 84:23]
  wire  _T_72 = block & dmaEn_0; // @[DMACtrlWRMask.scala 88:15]
  wire  _T_78 = 2'h1 == rState; // @[Mux.scala 80:60]
  wire  _T_80 = 2'h2 == rState; // @[Mux.scala 80:60]
  wire  _T_82 = 2'h3 == rState; // @[Mux.scala 80:60]
  wire  isReq = rState == 2'h1; // @[DMACtrlWRMask.scala 120:22]
  wire  isData = rState == 2'h2; // @[DMACtrlWRMask.scala 121:23]
  wire  isBlock = rState == 2'h3; // @[DMACtrlWRMask.scala 122:24]
  wire [63:0] _T_84 = dmaEn_0 ? dmaAXIAddr : {{32'd0}, dmaAXIAddrR}; // @[DMACtrlWRMask.scala 126:26]
  wire  _T_88 = isReq | isData; // @[DMACtrlWRMask.scala 132:30]
  reg [8:0] wCnt; // @[DMACtrlWRMask.scala 137:22]
  reg [2:0] wState; // @[DMACtrlWRMask.scala 139:23]
  wire  isWIdle = wState == 3'h0; // @[DMACtrlWRMask.scala 142:24]
  wire  isWReq = wState == 3'h1; // @[DMACtrlWRMask.scala 143:23]
  wire  isWData = wState == 3'h2; // @[DMACtrlWRMask.scala 144:24]
  wire  isWB = wState == 3'h3; // @[DMACtrlWRMask.scala 145:21]
  wire  isWBlock = wState == 3'h4; // @[DMACtrlWRMask.scala 146:25]
  wire  _T_90 = dmaEnWR_0 & changeState; // @[DMACtrlWRMask.scala 149:13]
  wire  _T_91 = io_dataIn_wready & io_dataIn_wlast; // @[DMACtrlWRMask.scala 154:47]
  wire  _T_92 = _T_91 & io_dataOutMMIO_ready; // @[DMACtrlWRMask.scala 154:66]
  wire [1:0] _T_93 = {io_dataIn_awready,_T_92}; // @[Cat.scala 29:58]
  wire  _T_94 = 2'h2 == _T_93; // @[Mux.scala 80:60]
  wire  _T_96 = 2'h3 == _T_93; // @[Mux.scala 80:60]
  wire  _T_100 = 3'h0 == wState; // @[Mux.scala 80:60]
  wire  _T_102 = 3'h1 == wState; // @[Mux.scala 80:60]
  wire  _T_104 = 3'h2 == wState; // @[Mux.scala 80:60]
  wire  _T_106 = 3'h3 == wState; // @[Mux.scala 80:60]
  wire  _T_108 = 3'h4 == wState; // @[Mux.scala 80:60]
  wire  _T_111 = isWData | isWReq; // @[DMACtrlWRMask.scala 201:40]
  wire  _T_112 = io_dataOutMMIO_ready & _T_111; // @[DMACtrlWRMask.scala 201:28]
  wire  _T_113 = _T_112 & io_dataIn_wready; // @[DMACtrlWRMask.scala 201:51]
  wire [8:0] _T_115 = wCnt + 9'h1; // @[DMACtrlWRMask.scala 202:12]
  wire [31:0] _GEN_0 = {{23'd0}, wCnt}; // @[DMACtrlWRMask.scala 212:27]
  wire  _T_121 = isWIdle & dmaEnWR_0; // @[DMACtrlWRMask.scala 217:38]
  wire  _T_122 = _T_121 & changeState; // @[DMACtrlWRMask.scala 217:49]
  wire  _T_127 = isWB & io_dataIn_bvalid; // @[DMACtrlWRMask.scala 225:12]
  wire  _T_130 = _T_88 & io_dataIn_rlast; // @[DMACtrlWRMask.scala 231:25]
  wire  _T_131 = _T_130 & dmaEnWR_0; // @[DMACtrlWRMask.scala 231:44]
  wire  _T_132 = _T_131 | changeState; // @[DMACtrlWRMask.scala 230:8]
  wire  _T_134 = ~io_dataIn_bvalid; // @[DMACtrlWRMask.scala 251:27]
  wire  _T_135 = dmaEnWR_0 & _T_134; // @[DMACtrlWRMask.scala 251:24]
  wire  _T_136 = ~isWBlock; // @[DMACtrlWRMask.scala 251:48]
  wire  _T_137 = _T_135 & _T_136; // @[DMACtrlWRMask.scala 251:45]
  wire  _T_138 = ~io_dataIn_rlast; // @[DMACtrlWRMask.scala 251:71]
  wire  _T_139 = dmaEn_0 & _T_138; // @[DMACtrlWRMask.scala 251:68]
  wire  _T_140 = ~isBlock; // @[DMACtrlWRMask.scala 251:91]
  wire  _T_141 = _T_139 & _T_140; // @[DMACtrlWRMask.scala 251:88]
  wire  _T_142 = _T_137 | _T_141; // @[DMACtrlWRMask.scala 251:58]
  wire  _T_144 = _T_88 | isWReq; // @[DMACtrlWRMask.scala 256:33]
  wire  _T_145 = _T_144 | isWData; // @[DMACtrlWRMask.scala 256:42]
  wire  DMABuzy = _T_145 | isWB; // @[DMACtrlWRMask.scala 256:53]
  wire  _T_146 = dmaEn_0 & isCfg; // @[DMACtrlWRMask.scala 277:35]
  wire  _T_147 = isWReq | isWData; // @[DMACtrlWRMask.scala 277:67]
  wire [31:0] CGRAOutAddr = portArbitInst_io_out; // @[DMACtrlWRMask.scala 54:25 DMACtrlWRMask.scala 63:15]
  wire [31:0] _T_148 = _T_147 ? CGRAOutAddr : 32'h2010000; // @[DMACtrlWRMask.scala 277:59]
  wire [63:0] _T_149 = _T_146 ? dmaDstAddr : {{32'd0}, _T_148}; // @[DMACtrlWRMask.scala 277:28]
  wire  _T_152 = _T_88 & io_dataIn_rvalid; // @[DMACtrlWRMask.scala 284:46]
  wire  blockDMA = _T_142; // @[DMACtrlWRMask.scala 250:22 DMACtrlWRMask.scala 251:12]
  adresPortArbit portArbitInst ( // @[DMACtrlWRMask.scala 56:29]
    .clock(portArbitInst_clock),
    .reset(portArbitInst_reset),
    .io_regEn(portArbitInst_io_regEn),
    .io_in_0_valid(portArbitInst_io_in_0_valid),
    .io_in_1_valid(portArbitInst_io_in_1_valid),
    .io_in_2_valid(portArbitInst_io_in_2_valid),
    .io_in_3_valid(portArbitInst_io_in_3_valid),
    .io_in_4_valid(portArbitInst_io_in_4_valid),
    .io_in_5_valid(portArbitInst_io_in_5_valid),
    .io_in_6_valid(portArbitInst_io_in_6_valid),
    .io_in_7_valid(portArbitInst_io_in_7_valid),
    .io_in_8_valid(portArbitInst_io_in_8_valid),
    .io_in_9_valid(portArbitInst_io_in_9_valid),
    .io_in_10_valid(portArbitInst_io_in_10_valid),
    .io_in_11_valid(portArbitInst_io_in_11_valid),
    .io_in_12_valid(portArbitInst_io_in_12_valid),
    .io_in_13_valid(portArbitInst_io_in_13_valid),
    .io_in_14_valid(portArbitInst_io_in_14_valid),
    .io_in_15_valid(portArbitInst_io_in_15_valid),
    .io_dmaEn(portArbitInst_io_dmaEn),
    .io_out(portArbitInst_io_out)
  );
  assign io_dataIn_awvalid = wState == 3'h1; // @[DMACtrlWRMask.scala 187:21]
  assign io_dataIn_awaddr = dmaCtrl_0[63:32]; // @[DMACtrlWRMask.scala 188:20]
  assign io_dataIn_awlen = dmaLenW[7:0]; // @[DMACtrlWRMask.scala 190:19]
  assign io_dataIn_wvalid = io_dataOutMMIO_ready & _T_111; // @[DMACtrlWRMask.scala 209:20]
  assign io_dataIn_wdata = io_dataOutMMIO_data_read; // @[DMACtrlWRMask.scala 210:19]
  assign io_dataIn_wlast = _GEN_0 == dmaLenW; // @[DMACtrlWRMask.scala 212:19]
  assign io_dataIn_bready = wState == 3'h3; // @[DMACtrlWRMask.scala 215:20]
  assign io_dataIn_arvalid = rState == 2'h1; // @[DMACtrlWRMask.scala 125:21]
  assign io_dataIn_araddr = _T_84[31:0]; // @[DMACtrlWRMask.scala 126:20]
  assign io_dataIn_arlen = dmaEn_0 ? dmaLen[7:0] : dmaLenR[7:0]; // @[DMACtrlWRMask.scala 128:19]
  assign io_dataIn_rready = _T_88 & io_dataOutMMIO_ready; // @[DMACtrlWRMask.scala 132:20]
  assign io_dataOutMMIO_valid = _T_152 | _T_147; // @[DMACtrlWRMask.scala 284:24]
  assign io_dataOutMMIO_data_write = io_dataIn_rdata; // @[DMACtrlWRMask.scala 286:29]
  assign io_dataOutMMIO_wen = isData & io_dataIn_rvalid; // @[DMACtrlWRMask.scala 279:22]
  assign io_dataOutMMIO_addr = _T_149[31:0]; // @[DMACtrlWRMask.scala 277:23]
  assign blockDMA_0 = blockDMA;
  assign DMABuzy_0 = DMABuzy;
  assign portArbitInst_clock = clock;
  assign portArbitInst_reset = reset;
  assign portArbitInst_io_regEn = _T_122 | _T_113; // @[DMACtrlWRMask.scala 217:26]
  assign portArbitInst_io_in_0_valid = dmaCGRAOutMask[0]; // @[DMACtrlWRMask.scala 59:34]
  assign portArbitInst_io_in_1_valid = dmaCGRAOutMask[1]; // @[DMACtrlWRMask.scala 59:34]
  assign portArbitInst_io_in_2_valid = dmaCGRAOutMask[2]; // @[DMACtrlWRMask.scala 59:34]
  assign portArbitInst_io_in_3_valid = dmaCGRAOutMask[3]; // @[DMACtrlWRMask.scala 59:34]
  assign portArbitInst_io_in_4_valid = dmaCGRAOutMask[4]; // @[DMACtrlWRMask.scala 59:34]
  assign portArbitInst_io_in_5_valid = dmaCGRAOutMask[5]; // @[DMACtrlWRMask.scala 59:34]
  assign portArbitInst_io_in_6_valid = dmaCGRAOutMask[6]; // @[DMACtrlWRMask.scala 59:34]
  assign portArbitInst_io_in_7_valid = dmaCGRAOutMask[7]; // @[DMACtrlWRMask.scala 59:34]
  assign portArbitInst_io_in_8_valid = dmaCGRAOutMask[8]; // @[DMACtrlWRMask.scala 59:34]
  assign portArbitInst_io_in_9_valid = dmaCGRAOutMask[9]; // @[DMACtrlWRMask.scala 59:34]
  assign portArbitInst_io_in_10_valid = dmaCGRAOutMask[10]; // @[DMACtrlWRMask.scala 59:34]
  assign portArbitInst_io_in_11_valid = dmaCGRAOutMask[11]; // @[DMACtrlWRMask.scala 59:34]
  assign portArbitInst_io_in_12_valid = dmaCGRAOutMask[12]; // @[DMACtrlWRMask.scala 59:34]
  assign portArbitInst_io_in_13_valid = dmaCGRAOutMask[13]; // @[DMACtrlWRMask.scala 59:34]
  assign portArbitInst_io_in_14_valid = dmaCGRAOutMask[14]; // @[DMACtrlWRMask.scala 59:34]
  assign portArbitInst_io_in_15_valid = dmaCGRAOutMask[15]; // @[DMACtrlWRMask.scala 59:34]
  assign portArbitInst_io_dmaEn = dmaEnWR_0; // @[DMACtrlWRMask.scala 62:26]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  changeState = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  rState = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  dmaNext = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  wCnt = _RAND_3[8:0];
  _RAND_4 = {1{`RANDOM}};
  wState = _RAND_4[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      changeState <= 1'h0;
    end else if (changeState) begin
      if (_T_127) begin
        changeState <= 1'h0;
      end
    end else begin
      changeState <= _T_132;
    end
    if (reset) begin
      rState <= 2'h0;
    end else if (_T_82) begin
      if (_T_72) begin
        rState <= 2'h3;
      end else begin
        rState <= 2'h0;
      end
    end else if (_T_80) begin
      if (io_dataIn_rlast) begin
        if (_T_72) begin
          rState <= 2'h3;
        end else begin
          rState <= 2'h0;
        end
      end else begin
        rState <= 2'h2;
      end
    end else if (_T_78) begin
      if (_T_71) begin
        if (io_dataIn_rlast) begin
          if (_T_72) begin
            rState <= 2'h3;
          end else begin
            rState <= 2'h0;
          end
        end else begin
          rState <= 2'h2;
        end
      end else begin
        rState <= 2'h1;
      end
    end else if (_T_69) begin
      rState <= 2'h1;
    end else begin
      rState <= 2'h0;
    end
    dmaNext <= dmaEn_0 | dmaEnWR_0;
    if (reset) begin
      wCnt <= 9'h0;
    end else if (isWIdle) begin
      wCnt <= 9'h0;
    end else if (_T_113) begin
      wCnt <= _T_115;
    end
    if (reset) begin
      wState <= 3'h0;
    end else if (_T_108) begin
      if (block) begin
        wState <= 3'h4;
      end else begin
        wState <= 3'h0;
      end
    end else if (_T_106) begin
      if (io_dataIn_bvalid) begin
        if (block) begin
          wState <= 3'h4;
        end else begin
          wState <= 3'h0;
        end
      end else begin
        wState <= 3'h3;
      end
    end else if (_T_104) begin
      if (_T_92) begin
        wState <= 3'h3;
      end else begin
        wState <= 3'h2;
      end
    end else if (_T_102) begin
      if (_T_96) begin
        wState <= 3'h3;
      end else if (_T_94) begin
        wState <= 3'h2;
      end else begin
        wState <= 3'h1;
      end
    end else if (_T_100) begin
      if (_T_90) begin
        wState <= 3'h1;
      end else begin
        wState <= 3'h0;
      end
    end
  end
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram [0:19]; // @[Decoupled.scala 209:16]
  wire [31:0] ram__T_11_data; // @[Decoupled.scala 209:16]
  wire [4:0] ram__T_11_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram__T_3_data; // @[Decoupled.scala 209:16]
  wire [4:0] ram__T_3_addr; // @[Decoupled.scala 209:16]
  wire  ram__T_3_mask; // @[Decoupled.scala 209:16]
  wire  ram__T_3_en; // @[Decoupled.scala 209:16]
  reg [4:0] enq_ptr_value; // @[Counter.scala 29:33]
  reg [4:0] deq_ptr_value; // @[Counter.scala 29:33]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 214:33]
  wire  _T = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  empty = ptr_match & _T; // @[Decoupled.scala 215:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 216:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  wrap = enq_ptr_value == 5'h13; // @[Counter.scala 38:24]
  wire [4:0] _T_5 = enq_ptr_value + 5'h1; // @[Counter.scala 39:22]
  wire  wrap_1 = deq_ptr_value == 5'h13; // @[Counter.scala 38:24]
  wire [4:0] _T_7 = deq_ptr_value + 5'h1; // @[Counter.scala 39:22]
  wire  _T_8 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  assign ram__T_11_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram__T_11_data = ram[ram__T_11_addr]; // @[Decoupled.scala 209:16]
  `else
  assign ram__T_11_data = ram__T_11_addr >= 5'h14 ? _RAND_1[31:0] : ram[ram__T_11_addr]; // @[Decoupled.scala 209:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram__T_3_data = io_enq_bits;
  assign ram__T_3_addr = enq_ptr_value;
  assign ram__T_3_mask = 1'h1;
  assign ram__T_3_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits = ram__T_11_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 20; initvar = initvar+1)
    ram[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enq_ptr_value = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  deq_ptr_value = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram__T_3_en & ram__T_3_mask) begin
      ram[ram__T_3_addr] <= ram__T_3_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      enq_ptr_value <= 5'h0;
    end else if (do_enq) begin
      if (wrap) begin
        enq_ptr_value <= 5'h0;
      end else begin
        enq_ptr_value <= _T_5;
      end
    end
    if (reset) begin
      deq_ptr_value <= 5'h0;
    end else if (do_deq) begin
      if (wrap_1) begin
        deq_ptr_value <= 5'h0;
      end else begin
        deq_ptr_value <= _T_7;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_8) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module adressGenIn(
  input        clock,
  input        reset,
  input        io_validList_0,
  input        io_validList_1,
  input        io_validList_2,
  input        io_validList_3,
  input        io_validList_4,
  input        io_validList_5,
  input        io_validList_6,
  input        io_validList_7,
  input        io_validList_8,
  input        io_validList_9,
  input        io_validList_10,
  input        io_validList_11,
  input        io_validList_12,
  input        io_validList_13,
  input        io_validList_14,
  input        io_update,
  input        io_clear,
  output [3:0] io_sel1,
  output [3:0] io_sel2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [3:0] _T = io_validList_14 ? 4'he : 4'hf; // @[Mux.scala 47:69]
  wire [3:0] _T_1 = io_validList_13 ? 4'hd : _T; // @[Mux.scala 47:69]
  wire [3:0] _T_2 = io_validList_12 ? 4'hc : _T_1; // @[Mux.scala 47:69]
  wire [3:0] _T_3 = io_validList_11 ? 4'hb : _T_2; // @[Mux.scala 47:69]
  wire [3:0] _T_4 = io_validList_10 ? 4'ha : _T_3; // @[Mux.scala 47:69]
  wire [3:0] _T_5 = io_validList_9 ? 4'h9 : _T_4; // @[Mux.scala 47:69]
  wire [3:0] _T_6 = io_validList_8 ? 4'h8 : _T_5; // @[Mux.scala 47:69]
  wire [3:0] _T_7 = io_validList_7 ? 4'h7 : _T_6; // @[Mux.scala 47:69]
  wire [3:0] _T_8 = io_validList_6 ? 4'h6 : _T_7; // @[Mux.scala 47:69]
  wire [3:0] _T_9 = io_validList_5 ? 4'h5 : _T_8; // @[Mux.scala 47:69]
  wire [3:0] _T_10 = io_validList_4 ? 4'h4 : _T_9; // @[Mux.scala 47:69]
  wire [3:0] _T_11 = io_validList_3 ? 4'h3 : _T_10; // @[Mux.scala 47:69]
  wire [3:0] _T_12 = io_validList_2 ? 4'h2 : _T_11; // @[Mux.scala 47:69]
  wire [3:0] _T_13 = io_validList_1 ? 4'h1 : _T_12; // @[Mux.scala 47:69]
  wire [3:0] _T_14 = io_validList_0 ? 4'h0 : _T_13; // @[Mux.scala 47:69]
  wire  _T_121 = io_clear | reset; // @[adressGenIn.scala 41:22]
  reg [3:0] indexSelReg; // @[Reg.scala 27:20]
  wire  _T_153 = 4'hf == indexSelReg; // @[Mux.scala 80:60]
  wire  _T_151 = 4'he == indexSelReg; // @[Mux.scala 80:60]
  wire  _T_149 = 4'hd == indexSelReg; // @[Mux.scala 80:60]
  wire  _T_147 = 4'hc == indexSelReg; // @[Mux.scala 80:60]
  wire  _T_145 = 4'hb == indexSelReg; // @[Mux.scala 80:60]
  wire  _T_143 = 4'ha == indexSelReg; // @[Mux.scala 80:60]
  wire  _T_141 = 4'h9 == indexSelReg; // @[Mux.scala 80:60]
  wire  _T_139 = 4'h8 == indexSelReg; // @[Mux.scala 80:60]
  wire  _T_137 = 4'h7 == indexSelReg; // @[Mux.scala 80:60]
  wire  _T_135 = 4'h6 == indexSelReg; // @[Mux.scala 80:60]
  wire  _T_133 = 4'h5 == indexSelReg; // @[Mux.scala 80:60]
  wire  _T_131 = 4'h4 == indexSelReg; // @[Mux.scala 80:60]
  wire  _T_129 = 4'h3 == indexSelReg; // @[Mux.scala 80:60]
  wire  _T_127 = 4'h2 == indexSelReg; // @[Mux.scala 80:60]
  wire  _T_125 = 4'h1 == indexSelReg; // @[Mux.scala 80:60]
  wire [3:0] _T_126 = _T_125 ? _T_13 : _T_14; // @[Mux.scala 80:57]
  wire [3:0] _T_128 = _T_127 ? _T_12 : _T_126; // @[Mux.scala 80:57]
  wire [3:0] _T_130 = _T_129 ? _T_11 : _T_128; // @[Mux.scala 80:57]
  wire [3:0] _T_132 = _T_131 ? _T_10 : _T_130; // @[Mux.scala 80:57]
  wire [3:0] _T_134 = _T_133 ? _T_9 : _T_132; // @[Mux.scala 80:57]
  wire [3:0] _T_136 = _T_135 ? _T_8 : _T_134; // @[Mux.scala 80:57]
  wire [3:0] _T_138 = _T_137 ? _T_7 : _T_136; // @[Mux.scala 80:57]
  wire [3:0] _T_140 = _T_139 ? _T_6 : _T_138; // @[Mux.scala 80:57]
  wire [3:0] _T_142 = _T_141 ? _T_5 : _T_140; // @[Mux.scala 80:57]
  wire [3:0] _T_144 = _T_143 ? _T_4 : _T_142; // @[Mux.scala 80:57]
  wire [3:0] _T_146 = _T_145 ? _T_3 : _T_144; // @[Mux.scala 80:57]
  wire [3:0] _T_148 = _T_147 ? _T_2 : _T_146; // @[Mux.scala 80:57]
  wire [3:0] _T_150 = _T_149 ? _T_1 : _T_148; // @[Mux.scala 80:57]
  wire [3:0] _T_152 = _T_151 ? _T : _T_150; // @[Mux.scala 80:57]
  wire [3:0] indexSelL = _T_153 ? 4'hf : _T_152; // @[Mux.scala 80:57]
  wire [3:0] _T_156 = indexSelL + 4'h1; // @[adressGenIn.scala 51:15]
  wire  _T_185 = 4'hf == _T_156; // @[Mux.scala 80:60]
  wire  _T_183 = 4'he == _T_156; // @[Mux.scala 80:60]
  wire  _T_181 = 4'hd == _T_156; // @[Mux.scala 80:60]
  wire  _T_179 = 4'hc == _T_156; // @[Mux.scala 80:60]
  wire  _T_177 = 4'hb == _T_156; // @[Mux.scala 80:60]
  wire  _T_175 = 4'ha == _T_156; // @[Mux.scala 80:60]
  wire  _T_173 = 4'h9 == _T_156; // @[Mux.scala 80:60]
  wire  _T_171 = 4'h8 == _T_156; // @[Mux.scala 80:60]
  wire  _T_169 = 4'h7 == _T_156; // @[Mux.scala 80:60]
  wire  _T_167 = 4'h6 == _T_156; // @[Mux.scala 80:60]
  wire  _T_165 = 4'h5 == _T_156; // @[Mux.scala 80:60]
  wire  _T_163 = 4'h4 == _T_156; // @[Mux.scala 80:60]
  wire  _T_161 = 4'h3 == _T_156; // @[Mux.scala 80:60]
  wire  _T_159 = 4'h2 == _T_156; // @[Mux.scala 80:60]
  wire  _T_157 = 4'h1 == _T_156; // @[Mux.scala 80:60]
  wire [3:0] _T_158 = _T_157 ? _T_13 : _T_14; // @[Mux.scala 80:57]
  wire [3:0] _T_160 = _T_159 ? _T_12 : _T_158; // @[Mux.scala 80:57]
  wire [3:0] _T_162 = _T_161 ? _T_11 : _T_160; // @[Mux.scala 80:57]
  wire [3:0] _T_164 = _T_163 ? _T_10 : _T_162; // @[Mux.scala 80:57]
  wire [3:0] _T_166 = _T_165 ? _T_9 : _T_164; // @[Mux.scala 80:57]
  wire [3:0] _T_168 = _T_167 ? _T_8 : _T_166; // @[Mux.scala 80:57]
  wire [3:0] _T_170 = _T_169 ? _T_7 : _T_168; // @[Mux.scala 80:57]
  wire [3:0] _T_172 = _T_171 ? _T_6 : _T_170; // @[Mux.scala 80:57]
  wire [3:0] _T_174 = _T_173 ? _T_5 : _T_172; // @[Mux.scala 80:57]
  wire [3:0] _T_176 = _T_175 ? _T_4 : _T_174; // @[Mux.scala 80:57]
  wire [3:0] _T_178 = _T_177 ? _T_3 : _T_176; // @[Mux.scala 80:57]
  wire [3:0] _T_180 = _T_179 ? _T_2 : _T_178; // @[Mux.scala 80:57]
  wire [3:0] _T_182 = _T_181 ? _T_1 : _T_180; // @[Mux.scala 80:57]
  wire [3:0] _T_184 = _T_183 ? _T : _T_182; // @[Mux.scala 80:57]
  wire [3:0] indexSelH = _T_185 ? 4'hf : _T_184; // @[Mux.scala 80:57]
  wire [3:0] _T_123 = indexSelH + 4'h1; // @[adressGenIn.scala 42:40]
  assign io_sel1 = _T_153 ? 4'hf : _T_152; // @[adressGenIn.scala 56:11]
  assign io_sel2 = _T_185 ? 4'hf : _T_184; // @[adressGenIn.scala 57:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  indexSelReg = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_121) begin
      indexSelReg <= 4'h0;
    end else if (io_update) begin
      indexSelReg <= _T_123;
    end
  end
endmodule
module SynInMask(
  input          clock,
  input          reset,
  input          io_valid,
  output         io_ready,
  input  [63:0]  io_dataIn,
  output [32:0]  io_dataOut_0,
  output [32:0]  io_dataOut_1,
  output [32:0]  io_dataOut_2,
  output [32:0]  io_dataOut_3,
  output [32:0]  io_dataOut_4,
  output [32:0]  io_dataOut_5,
  output [32:0]  io_dataOut_6,
  output [32:0]  io_dataOut_7,
  output [32:0]  io_dataOut_8,
  output [32:0]  io_dataOut_9,
  output [32:0]  io_dataOut_10,
  output [32:0]  io_dataOut_11,
  output [32:0]  io_dataOut_12,
  output [32:0]  io_dataOut_13,
  output [32:0]  io_dataOut_14,
  output [32:0]  io_dataOut_15,
  input          io_delayen,
  input  [63:0]  io_delayCycle,
  input          dmaEnWR_0,
  input  [191:0] dmaCtrl_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
`endif // RANDOMIZE_REG_INIT
  wire  adrGenInst_clock; // @[SynInMask.scala 28:25]
  wire  adrGenInst_reset; // @[SynInMask.scala 28:25]
  wire  adrGenInst_io_validList_0; // @[SynInMask.scala 28:25]
  wire  adrGenInst_io_validList_1; // @[SynInMask.scala 28:25]
  wire  adrGenInst_io_validList_2; // @[SynInMask.scala 28:25]
  wire  adrGenInst_io_validList_3; // @[SynInMask.scala 28:25]
  wire  adrGenInst_io_validList_4; // @[SynInMask.scala 28:25]
  wire  adrGenInst_io_validList_5; // @[SynInMask.scala 28:25]
  wire  adrGenInst_io_validList_6; // @[SynInMask.scala 28:25]
  wire  adrGenInst_io_validList_7; // @[SynInMask.scala 28:25]
  wire  adrGenInst_io_validList_8; // @[SynInMask.scala 28:25]
  wire  adrGenInst_io_validList_9; // @[SynInMask.scala 28:25]
  wire  adrGenInst_io_validList_10; // @[SynInMask.scala 28:25]
  wire  adrGenInst_io_validList_11; // @[SynInMask.scala 28:25]
  wire  adrGenInst_io_validList_12; // @[SynInMask.scala 28:25]
  wire  adrGenInst_io_validList_13; // @[SynInMask.scala 28:25]
  wire  adrGenInst_io_validList_14; // @[SynInMask.scala 28:25]
  wire  adrGenInst_io_update; // @[SynInMask.scala 28:25]
  wire  adrGenInst_io_clear; // @[SynInMask.scala 28:25]
  wire [3:0] adrGenInst_io_sel1; // @[SynInMask.scala 28:25]
  wire [3:0] adrGenInst_io_sel2; // @[SynInMask.scala 28:25]
  wire  dmaCGRAInMask_0 = dmaCtrl_0[64]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_1 = dmaCtrl_0[65]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_2 = dmaCtrl_0[66]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_3 = dmaCtrl_0[67]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_4 = dmaCtrl_0[68]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_5 = dmaCtrl_0[69]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_6 = dmaCtrl_0[70]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_7 = dmaCtrl_0[71]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_8 = dmaCtrl_0[72]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_9 = dmaCtrl_0[73]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_10 = dmaCtrl_0[74]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_11 = dmaCtrl_0[75]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_12 = dmaCtrl_0[76]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_13 = dmaCtrl_0[77]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_14 = dmaCtrl_0[78]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_15 = dmaCtrl_0[79]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_16 = dmaCtrl_0[80]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_17 = dmaCtrl_0[81]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_18 = dmaCtrl_0[82]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_19 = dmaCtrl_0[83]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_20 = dmaCtrl_0[84]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_21 = dmaCtrl_0[85]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_22 = dmaCtrl_0[86]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_23 = dmaCtrl_0[87]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_24 = dmaCtrl_0[88]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_25 = dmaCtrl_0[89]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_26 = dmaCtrl_0[90]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_27 = dmaCtrl_0[91]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_28 = dmaCtrl_0[92]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_29 = dmaCtrl_0[93]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_30 = dmaCtrl_0[94]; // @[SynInMask.scala 30:59]
  wire  dmaCGRAInMask_31 = dmaCtrl_0[95]; // @[SynInMask.scala 30:59]
  wire [5:0] _T_1 = {{5'd0}, dmaCGRAInMask_0}; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_35 = {{4'd0}, dmaCGRAInMask_1}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_4 = _T_1[4:0] + _GEN_35; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_36 = {{4'd0}, dmaCGRAInMask_2}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_6 = _T_4 + _GEN_36; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_37 = {{4'd0}, dmaCGRAInMask_3}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_8 = _T_6 + _GEN_37; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_38 = {{4'd0}, dmaCGRAInMask_4}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_10 = _T_8 + _GEN_38; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_39 = {{4'd0}, dmaCGRAInMask_5}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_12 = _T_10 + _GEN_39; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_40 = {{4'd0}, dmaCGRAInMask_6}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_14 = _T_12 + _GEN_40; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_41 = {{4'd0}, dmaCGRAInMask_7}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_16 = _T_14 + _GEN_41; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_42 = {{4'd0}, dmaCGRAInMask_8}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_18 = _T_16 + _GEN_42; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_43 = {{4'd0}, dmaCGRAInMask_9}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_20 = _T_18 + _GEN_43; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_44 = {{4'd0}, dmaCGRAInMask_10}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_22 = _T_20 + _GEN_44; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_45 = {{4'd0}, dmaCGRAInMask_11}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_24 = _T_22 + _GEN_45; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_46 = {{4'd0}, dmaCGRAInMask_12}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_26 = _T_24 + _GEN_46; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_47 = {{4'd0}, dmaCGRAInMask_13}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_28 = _T_26 + _GEN_47; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_48 = {{4'd0}, dmaCGRAInMask_14}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_30 = _T_28 + _GEN_48; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_49 = {{4'd0}, dmaCGRAInMask_15}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_32 = _T_30 + _GEN_49; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_50 = {{4'd0}, dmaCGRAInMask_16}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_34 = _T_32 + _GEN_50; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_51 = {{4'd0}, dmaCGRAInMask_17}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_36 = _T_34 + _GEN_51; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_52 = {{4'd0}, dmaCGRAInMask_18}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_38 = _T_36 + _GEN_52; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_53 = {{4'd0}, dmaCGRAInMask_19}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_40 = _T_38 + _GEN_53; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_54 = {{4'd0}, dmaCGRAInMask_20}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_42 = _T_40 + _GEN_54; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_55 = {{4'd0}, dmaCGRAInMask_21}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_44 = _T_42 + _GEN_55; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_56 = {{4'd0}, dmaCGRAInMask_22}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_46 = _T_44 + _GEN_56; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_57 = {{4'd0}, dmaCGRAInMask_23}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_48 = _T_46 + _GEN_57; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_58 = {{4'd0}, dmaCGRAInMask_24}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_50 = _T_48 + _GEN_58; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_59 = {{4'd0}, dmaCGRAInMask_25}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_52 = _T_50 + _GEN_59; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_60 = {{4'd0}, dmaCGRAInMask_26}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_54 = _T_52 + _GEN_60; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_61 = {{4'd0}, dmaCGRAInMask_27}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_56 = _T_54 + _GEN_61; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_62 = {{4'd0}, dmaCGRAInMask_28}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_58 = _T_56 + _GEN_62; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_63 = {{4'd0}, dmaCGRAInMask_29}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_60 = _T_58 + _GEN_63; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_64 = {{4'd0}, dmaCGRAInMask_30}; // @[SynInMask.scala 33:58]
  wire [4:0] _T_62 = _T_60 + _GEN_64; // @[SynInMask.scala 33:58]
  wire [4:0] _GEN_65 = {{4'd0}, dmaCGRAInMask_31}; // @[SynInMask.scala 33:58]
  wire [4:0] ones = _T_62 + _GEN_65; // @[SynInMask.scala 33:58]
  wire [3:0] _T_68 = ones[4:1] + 4'h1; // @[SynInMask.scala 34:51]
  wire [3:0] clearCount = ones[0] ? _T_68 : ones[4:1]; // @[SynInMask.scala 34:23]
  reg [3:0] clearCountReg; // @[Reg.scala 27:20]
  wire [3:0] _T_71 = clearCountReg + 4'h1; // @[SynInMask.scala 38:31]
  wire  clearUp = _T_71 == clearCount; // @[SynInMask.scala 38:37]
  wire  _T_678 = 4'hf == adrGenInst_io_sel1; // @[Mux.scala 80:60]
  reg  outValidsWire_15; // @[Reg.scala 27:20]
  wire  _T_630 = ~outValidsWire_15; // @[SynInMask.scala 84:25]
  wire  _T_618 = 4'hf == adrGenInst_io_sel2; // @[SynInMask.scala 80:22]
  wire  lastNoValid = ones[0] & clearUp; // @[SynInMask.scala 52:29]
  wire  _T_619 = ~lastNoValid; // @[SynInMask.scala 80:48]
  wire  _T_620 = _T_618 & _T_619; // @[SynInMask.scala 80:45]
  wire  _T_624 = _T_678 | _T_620; // @[SynInMask.scala 82:31]
  reg  outValidsWire_0; // @[Reg.scala 27:20]
  wire  _T_81 = ~dmaCGRAInMask_0; // @[SynInMask.scala 57:77]
  wire  rstList_0 = outValidsWire_0 | _T_81; // @[SynInMask.scala 57:73]
  reg  outValidsWire_1; // @[Reg.scala 27:20]
  wire  _T_82 = ~dmaCGRAInMask_1; // @[SynInMask.scala 57:77]
  wire  rstList_1 = outValidsWire_1 | _T_82; // @[SynInMask.scala 57:73]
  wire  _T_98 = rstList_0 & rstList_1; // @[SynInMask.scala 58:53]
  reg  outValidsWire_2; // @[Reg.scala 27:20]
  wire  _T_83 = ~dmaCGRAInMask_2; // @[SynInMask.scala 57:77]
  wire  rstList_2 = outValidsWire_2 | _T_83; // @[SynInMask.scala 57:73]
  wire  _T_99 = _T_98 & rstList_2; // @[SynInMask.scala 58:53]
  reg  outValidsWire_3; // @[Reg.scala 27:20]
  wire  _T_84 = ~dmaCGRAInMask_3; // @[SynInMask.scala 57:77]
  wire  rstList_3 = outValidsWire_3 | _T_84; // @[SynInMask.scala 57:73]
  wire  _T_100 = _T_99 & rstList_3; // @[SynInMask.scala 58:53]
  reg  outValidsWire_4; // @[Reg.scala 27:20]
  wire  _T_85 = ~dmaCGRAInMask_4; // @[SynInMask.scala 57:77]
  wire  rstList_4 = outValidsWire_4 | _T_85; // @[SynInMask.scala 57:73]
  wire  _T_101 = _T_100 & rstList_4; // @[SynInMask.scala 58:53]
  reg  outValidsWire_5; // @[Reg.scala 27:20]
  wire  _T_86 = ~dmaCGRAInMask_5; // @[SynInMask.scala 57:77]
  wire  rstList_5 = outValidsWire_5 | _T_86; // @[SynInMask.scala 57:73]
  wire  _T_102 = _T_101 & rstList_5; // @[SynInMask.scala 58:53]
  reg  outValidsWire_6; // @[Reg.scala 27:20]
  wire  _T_87 = ~dmaCGRAInMask_6; // @[SynInMask.scala 57:77]
  wire  rstList_6 = outValidsWire_6 | _T_87; // @[SynInMask.scala 57:73]
  wire  _T_103 = _T_102 & rstList_6; // @[SynInMask.scala 58:53]
  reg  outValidsWire_7; // @[Reg.scala 27:20]
  wire  _T_88 = ~dmaCGRAInMask_7; // @[SynInMask.scala 57:77]
  wire  rstList_7 = outValidsWire_7 | _T_88; // @[SynInMask.scala 57:73]
  wire  _T_104 = _T_103 & rstList_7; // @[SynInMask.scala 58:53]
  reg  outValidsWire_8; // @[Reg.scala 27:20]
  wire  _T_89 = ~dmaCGRAInMask_8; // @[SynInMask.scala 57:77]
  wire  rstList_8 = outValidsWire_8 | _T_89; // @[SynInMask.scala 57:73]
  wire  _T_105 = _T_104 & rstList_8; // @[SynInMask.scala 58:53]
  reg  outValidsWire_9; // @[Reg.scala 27:20]
  wire  _T_90 = ~dmaCGRAInMask_9; // @[SynInMask.scala 57:77]
  wire  rstList_9 = outValidsWire_9 | _T_90; // @[SynInMask.scala 57:73]
  wire  _T_106 = _T_105 & rstList_9; // @[SynInMask.scala 58:53]
  reg  outValidsWire_10; // @[Reg.scala 27:20]
  wire  _T_91 = ~dmaCGRAInMask_10; // @[SynInMask.scala 57:77]
  wire  rstList_10 = outValidsWire_10 | _T_91; // @[SynInMask.scala 57:73]
  wire  _T_107 = _T_106 & rstList_10; // @[SynInMask.scala 58:53]
  reg  outValidsWire_11; // @[Reg.scala 27:20]
  wire  _T_92 = ~dmaCGRAInMask_11; // @[SynInMask.scala 57:77]
  wire  rstList_11 = outValidsWire_11 | _T_92; // @[SynInMask.scala 57:73]
  wire  _T_108 = _T_107 & rstList_11; // @[SynInMask.scala 58:53]
  reg  outValidsWire_12; // @[Reg.scala 27:20]
  wire  _T_93 = ~dmaCGRAInMask_12; // @[SynInMask.scala 57:77]
  wire  rstList_12 = outValidsWire_12 | _T_93; // @[SynInMask.scala 57:73]
  wire  _T_109 = _T_108 & rstList_12; // @[SynInMask.scala 58:53]
  reg  outValidsWire_13; // @[Reg.scala 27:20]
  wire  _T_94 = ~dmaCGRAInMask_13; // @[SynInMask.scala 57:77]
  wire  rstList_13 = outValidsWire_13 | _T_94; // @[SynInMask.scala 57:73]
  wire  _T_110 = _T_109 & rstList_13; // @[SynInMask.scala 58:53]
  reg  outValidsWire_14; // @[Reg.scala 27:20]
  wire  _T_95 = ~dmaCGRAInMask_14; // @[SynInMask.scala 57:77]
  wire  rstList_14 = outValidsWire_14 | _T_95; // @[SynInMask.scala 57:73]
  wire  _T_111 = _T_110 & rstList_14; // @[SynInMask.scala 58:53]
  wire  _T_96 = ~dmaCGRAInMask_15; // @[SynInMask.scala 57:77]
  wire  rstList_15 = outValidsWire_15 | _T_96; // @[SynInMask.scala 57:73]
  wire  dataRst = _T_111 & rstList_15; // @[SynInMask.scala 58:53]
  wire  _T_625 = _T_624 & dataRst; // @[SynInMask.scala 82:41]
  wire  _T_631 = _T_630 | _T_625; // @[SynInMask.scala 84:42]
  reg [5:0] delayCnt; // @[Reg.scala 27:20]
  wire  noWait = delayCnt == 6'h0; // @[SynInMask.scala 72:25]
  wire  _T_632 = _T_631 & noWait; // @[SynInMask.scala 84:58]
  wire  readyList_15 = _T_632 & dmaCGRAInMask_15; // @[SynInMask.scala 84:68]
  wire  _T_676 = 4'he == adrGenInst_io_sel1; // @[Mux.scala 80:60]
  wire  _T_597 = ~outValidsWire_14; // @[SynInMask.scala 84:25]
  wire  _T_585 = 4'he == adrGenInst_io_sel2; // @[SynInMask.scala 80:22]
  wire  _T_587 = _T_585 & _T_619; // @[SynInMask.scala 80:45]
  wire  _T_591 = _T_676 | _T_587; // @[SynInMask.scala 82:31]
  wire  _T_592 = _T_591 & dataRst; // @[SynInMask.scala 82:41]
  wire  _T_598 = _T_597 | _T_592; // @[SynInMask.scala 84:42]
  wire  _T_599 = _T_598 & noWait; // @[SynInMask.scala 84:58]
  wire  readyList_14 = _T_599 & dmaCGRAInMask_14; // @[SynInMask.scala 84:68]
  wire  _T_674 = 4'hd == adrGenInst_io_sel1; // @[Mux.scala 80:60]
  wire  _T_564 = ~outValidsWire_13; // @[SynInMask.scala 84:25]
  wire  _T_552 = 4'hd == adrGenInst_io_sel2; // @[SynInMask.scala 80:22]
  wire  _T_554 = _T_552 & _T_619; // @[SynInMask.scala 80:45]
  wire  _T_558 = _T_674 | _T_554; // @[SynInMask.scala 82:31]
  wire  _T_559 = _T_558 & dataRst; // @[SynInMask.scala 82:41]
  wire  _T_565 = _T_564 | _T_559; // @[SynInMask.scala 84:42]
  wire  _T_566 = _T_565 & noWait; // @[SynInMask.scala 84:58]
  wire  readyList_13 = _T_566 & dmaCGRAInMask_13; // @[SynInMask.scala 84:68]
  wire  _T_672 = 4'hc == adrGenInst_io_sel1; // @[Mux.scala 80:60]
  wire  _T_531 = ~outValidsWire_12; // @[SynInMask.scala 84:25]
  wire  _T_519 = 4'hc == adrGenInst_io_sel2; // @[SynInMask.scala 80:22]
  wire  _T_521 = _T_519 & _T_619; // @[SynInMask.scala 80:45]
  wire  _T_525 = _T_672 | _T_521; // @[SynInMask.scala 82:31]
  wire  _T_526 = _T_525 & dataRst; // @[SynInMask.scala 82:41]
  wire  _T_532 = _T_531 | _T_526; // @[SynInMask.scala 84:42]
  wire  _T_533 = _T_532 & noWait; // @[SynInMask.scala 84:58]
  wire  readyList_12 = _T_533 & dmaCGRAInMask_12; // @[SynInMask.scala 84:68]
  wire  _T_670 = 4'hb == adrGenInst_io_sel1; // @[Mux.scala 80:60]
  wire  _T_498 = ~outValidsWire_11; // @[SynInMask.scala 84:25]
  wire  _T_486 = 4'hb == adrGenInst_io_sel2; // @[SynInMask.scala 80:22]
  wire  _T_488 = _T_486 & _T_619; // @[SynInMask.scala 80:45]
  wire  _T_492 = _T_670 | _T_488; // @[SynInMask.scala 82:31]
  wire  _T_493 = _T_492 & dataRst; // @[SynInMask.scala 82:41]
  wire  _T_499 = _T_498 | _T_493; // @[SynInMask.scala 84:42]
  wire  _T_500 = _T_499 & noWait; // @[SynInMask.scala 84:58]
  wire  readyList_11 = _T_500 & dmaCGRAInMask_11; // @[SynInMask.scala 84:68]
  wire  _T_668 = 4'ha == adrGenInst_io_sel1; // @[Mux.scala 80:60]
  wire  _T_465 = ~outValidsWire_10; // @[SynInMask.scala 84:25]
  wire  _T_453 = 4'ha == adrGenInst_io_sel2; // @[SynInMask.scala 80:22]
  wire  _T_455 = _T_453 & _T_619; // @[SynInMask.scala 80:45]
  wire  _T_459 = _T_668 | _T_455; // @[SynInMask.scala 82:31]
  wire  _T_460 = _T_459 & dataRst; // @[SynInMask.scala 82:41]
  wire  _T_466 = _T_465 | _T_460; // @[SynInMask.scala 84:42]
  wire  _T_467 = _T_466 & noWait; // @[SynInMask.scala 84:58]
  wire  readyList_10 = _T_467 & dmaCGRAInMask_10; // @[SynInMask.scala 84:68]
  wire  _T_666 = 4'h9 == adrGenInst_io_sel1; // @[Mux.scala 80:60]
  wire  _T_432 = ~outValidsWire_9; // @[SynInMask.scala 84:25]
  wire  _T_420 = 4'h9 == adrGenInst_io_sel2; // @[SynInMask.scala 80:22]
  wire  _T_422 = _T_420 & _T_619; // @[SynInMask.scala 80:45]
  wire  _T_426 = _T_666 | _T_422; // @[SynInMask.scala 82:31]
  wire  _T_427 = _T_426 & dataRst; // @[SynInMask.scala 82:41]
  wire  _T_433 = _T_432 | _T_427; // @[SynInMask.scala 84:42]
  wire  _T_434 = _T_433 & noWait; // @[SynInMask.scala 84:58]
  wire  readyList_9 = _T_434 & dmaCGRAInMask_9; // @[SynInMask.scala 84:68]
  wire  _T_664 = 4'h8 == adrGenInst_io_sel1; // @[Mux.scala 80:60]
  wire  _T_399 = ~outValidsWire_8; // @[SynInMask.scala 84:25]
  wire  _T_387 = 4'h8 == adrGenInst_io_sel2; // @[SynInMask.scala 80:22]
  wire  _T_389 = _T_387 & _T_619; // @[SynInMask.scala 80:45]
  wire  _T_393 = _T_664 | _T_389; // @[SynInMask.scala 82:31]
  wire  _T_394 = _T_393 & dataRst; // @[SynInMask.scala 82:41]
  wire  _T_400 = _T_399 | _T_394; // @[SynInMask.scala 84:42]
  wire  _T_401 = _T_400 & noWait; // @[SynInMask.scala 84:58]
  wire  readyList_8 = _T_401 & dmaCGRAInMask_8; // @[SynInMask.scala 84:68]
  wire  _T_662 = 4'h7 == adrGenInst_io_sel1; // @[Mux.scala 80:60]
  wire  _T_366 = ~outValidsWire_7; // @[SynInMask.scala 84:25]
  wire  _T_354 = 4'h7 == adrGenInst_io_sel2; // @[SynInMask.scala 80:22]
  wire  _T_356 = _T_354 & _T_619; // @[SynInMask.scala 80:45]
  wire  _T_360 = _T_662 | _T_356; // @[SynInMask.scala 82:31]
  wire  _T_361 = _T_360 & dataRst; // @[SynInMask.scala 82:41]
  wire  _T_367 = _T_366 | _T_361; // @[SynInMask.scala 84:42]
  wire  _T_368 = _T_367 & noWait; // @[SynInMask.scala 84:58]
  wire  readyList_7 = _T_368 & dmaCGRAInMask_7; // @[SynInMask.scala 84:68]
  wire  _T_660 = 4'h6 == adrGenInst_io_sel1; // @[Mux.scala 80:60]
  wire  _T_333 = ~outValidsWire_6; // @[SynInMask.scala 84:25]
  wire  _T_321 = 4'h6 == adrGenInst_io_sel2; // @[SynInMask.scala 80:22]
  wire  _T_323 = _T_321 & _T_619; // @[SynInMask.scala 80:45]
  wire  _T_327 = _T_660 | _T_323; // @[SynInMask.scala 82:31]
  wire  _T_328 = _T_327 & dataRst; // @[SynInMask.scala 82:41]
  wire  _T_334 = _T_333 | _T_328; // @[SynInMask.scala 84:42]
  wire  _T_335 = _T_334 & noWait; // @[SynInMask.scala 84:58]
  wire  readyList_6 = _T_335 & dmaCGRAInMask_6; // @[SynInMask.scala 84:68]
  wire  _T_658 = 4'h5 == adrGenInst_io_sel1; // @[Mux.scala 80:60]
  wire  _T_300 = ~outValidsWire_5; // @[SynInMask.scala 84:25]
  wire  _T_288 = 4'h5 == adrGenInst_io_sel2; // @[SynInMask.scala 80:22]
  wire  _T_290 = _T_288 & _T_619; // @[SynInMask.scala 80:45]
  wire  _T_294 = _T_658 | _T_290; // @[SynInMask.scala 82:31]
  wire  _T_295 = _T_294 & dataRst; // @[SynInMask.scala 82:41]
  wire  _T_301 = _T_300 | _T_295; // @[SynInMask.scala 84:42]
  wire  _T_302 = _T_301 & noWait; // @[SynInMask.scala 84:58]
  wire  readyList_5 = _T_302 & dmaCGRAInMask_5; // @[SynInMask.scala 84:68]
  wire  _T_656 = 4'h4 == adrGenInst_io_sel1; // @[Mux.scala 80:60]
  wire  _T_267 = ~outValidsWire_4; // @[SynInMask.scala 84:25]
  wire  _T_255 = 4'h4 == adrGenInst_io_sel2; // @[SynInMask.scala 80:22]
  wire  _T_257 = _T_255 & _T_619; // @[SynInMask.scala 80:45]
  wire  _T_261 = _T_656 | _T_257; // @[SynInMask.scala 82:31]
  wire  _T_262 = _T_261 & dataRst; // @[SynInMask.scala 82:41]
  wire  _T_268 = _T_267 | _T_262; // @[SynInMask.scala 84:42]
  wire  _T_269 = _T_268 & noWait; // @[SynInMask.scala 84:58]
  wire  readyList_4 = _T_269 & dmaCGRAInMask_4; // @[SynInMask.scala 84:68]
  wire  _T_654 = 4'h3 == adrGenInst_io_sel1; // @[Mux.scala 80:60]
  wire  _T_234 = ~outValidsWire_3; // @[SynInMask.scala 84:25]
  wire  _T_222 = 4'h3 == adrGenInst_io_sel2; // @[SynInMask.scala 80:22]
  wire  _T_224 = _T_222 & _T_619; // @[SynInMask.scala 80:45]
  wire  _T_228 = _T_654 | _T_224; // @[SynInMask.scala 82:31]
  wire  _T_229 = _T_228 & dataRst; // @[SynInMask.scala 82:41]
  wire  _T_235 = _T_234 | _T_229; // @[SynInMask.scala 84:42]
  wire  _T_236 = _T_235 & noWait; // @[SynInMask.scala 84:58]
  wire  readyList_3 = _T_236 & dmaCGRAInMask_3; // @[SynInMask.scala 84:68]
  wire  _T_652 = 4'h2 == adrGenInst_io_sel1; // @[Mux.scala 80:60]
  wire  _T_201 = ~outValidsWire_2; // @[SynInMask.scala 84:25]
  wire  _T_189 = 4'h2 == adrGenInst_io_sel2; // @[SynInMask.scala 80:22]
  wire  _T_191 = _T_189 & _T_619; // @[SynInMask.scala 80:45]
  wire  _T_195 = _T_652 | _T_191; // @[SynInMask.scala 82:31]
  wire  _T_196 = _T_195 & dataRst; // @[SynInMask.scala 82:41]
  wire  _T_202 = _T_201 | _T_196; // @[SynInMask.scala 84:42]
  wire  _T_203 = _T_202 & noWait; // @[SynInMask.scala 84:58]
  wire  readyList_2 = _T_203 & dmaCGRAInMask_2; // @[SynInMask.scala 84:68]
  wire  _T_650 = 4'h1 == adrGenInst_io_sel1; // @[Mux.scala 80:60]
  wire  _T_168 = ~outValidsWire_1; // @[SynInMask.scala 84:25]
  wire  _T_156 = 4'h1 == adrGenInst_io_sel2; // @[SynInMask.scala 80:22]
  wire  _T_158 = _T_156 & _T_619; // @[SynInMask.scala 80:45]
  wire  _T_162 = _T_650 | _T_158; // @[SynInMask.scala 82:31]
  wire  _T_163 = _T_162 & dataRst; // @[SynInMask.scala 82:41]
  wire  _T_169 = _T_168 | _T_163; // @[SynInMask.scala 84:42]
  wire  _T_170 = _T_169 & noWait; // @[SynInMask.scala 84:58]
  wire  readyList_1 = _T_170 & dmaCGRAInMask_1; // @[SynInMask.scala 84:68]
  wire  _T_135 = ~outValidsWire_0; // @[SynInMask.scala 84:25]
  wire  _T_122 = 4'h0 == adrGenInst_io_sel1; // @[SynInMask.scala 79:22]
  wire  _T_123 = 4'h0 == adrGenInst_io_sel2; // @[SynInMask.scala 80:22]
  wire  _T_125 = _T_123 & _T_619; // @[SynInMask.scala 80:45]
  wire  _T_129 = _T_122 | _T_125; // @[SynInMask.scala 82:31]
  wire  _T_130 = _T_129 & dataRst; // @[SynInMask.scala 82:41]
  wire  _T_136 = _T_135 | _T_130; // @[SynInMask.scala 84:42]
  wire  _T_137 = _T_136 & noWait; // @[SynInMask.scala 84:58]
  wire  readyList_0 = _T_137 & dmaCGRAInMask_0; // @[SynInMask.scala 84:68]
  wire  _T_651 = _T_650 ? readyList_1 : readyList_0; // @[Mux.scala 80:57]
  wire  _T_653 = _T_652 ? readyList_2 : _T_651; // @[Mux.scala 80:57]
  wire  _T_655 = _T_654 ? readyList_3 : _T_653; // @[Mux.scala 80:57]
  wire  _T_657 = _T_656 ? readyList_4 : _T_655; // @[Mux.scala 80:57]
  wire  _T_659 = _T_658 ? readyList_5 : _T_657; // @[Mux.scala 80:57]
  wire  _T_661 = _T_660 ? readyList_6 : _T_659; // @[Mux.scala 80:57]
  wire  _T_663 = _T_662 ? readyList_7 : _T_661; // @[Mux.scala 80:57]
  wire  _T_665 = _T_664 ? readyList_8 : _T_663; // @[Mux.scala 80:57]
  wire  _T_667 = _T_666 ? readyList_9 : _T_665; // @[Mux.scala 80:57]
  wire  _T_669 = _T_668 ? readyList_10 : _T_667; // @[Mux.scala 80:57]
  wire  _T_671 = _T_670 ? readyList_11 : _T_669; // @[Mux.scala 80:57]
  wire  _T_673 = _T_672 ? readyList_12 : _T_671; // @[Mux.scala 80:57]
  wire  _T_675 = _T_674 ? readyList_13 : _T_673; // @[Mux.scala 80:57]
  wire  _T_677 = _T_676 ? readyList_14 : _T_675; // @[Mux.scala 80:57]
  wire  readySel = _T_678 ? readyList_15 : _T_677; // @[Mux.scala 80:57]
  wire  updateWire = readySel & io_valid; // @[SynInMask.scala 98:25]
  reg [5:0] delayReg; // @[Reg.scala 27:20]
  wire  _T_113 = delayCnt != 6'h0; // @[SynInMask.scala 65:28]
  wire  _T_114 = dataRst | _T_113; // @[SynInMask.scala 65:16]
  wire  _T_115 = delayReg != delayCnt; // @[SynInMask.scala 65:49]
  wire  _T_116 = _T_114 & _T_115; // @[SynInMask.scala 65:37]
  wire [5:0] _T_118 = delayCnt + 6'h1; // @[SynInMask.scala 66:16]
  wire  _T_120 = delayReg != 6'h0; // @[SynInMask.scala 70:14]
  wire  _T_131 = ~_T_130; // @[SynInMask.scala 83:27]
  wire  _T_132 = dataRst & _T_131; // @[SynInMask.scala 83:24]
  wire  _T_134 = _T_132 | reset; // @[SynInMask.scala 83:42]
  wire  _T_141 = io_valid & _T_136; // @[SynInMask.scala 85:55]
  wire  _T_142 = _T_141 & noWait; // @[SynInMask.scala 85:92]
  wire  _T_144 = _T_142 & _T_129; // @[SynInMask.scala 85:102]
  wire  _T_145 = _T_144 & dmaCGRAInMask_0; // @[SynInMask.scala 85:122]
  reg [31:0] inDatasWire_0; // @[Reg.scala 27:20]
  wire  _T_149 = _T_136 & io_valid; // @[SynInMask.scala 86:90]
  wire  _T_150 = _T_149 & noWait; // @[SynInMask.scala 86:102]
  wire  _T_152 = _T_150 & _T_129; // @[SynInMask.scala 86:111]
  wire  _T_153 = _T_152 & dmaCGRAInMask_0; // @[SynInMask.scala 86:131]
  wire  _T_164 = ~_T_163; // @[SynInMask.scala 83:27]
  wire  _T_165 = dataRst & _T_164; // @[SynInMask.scala 83:24]
  wire  _T_167 = _T_165 | reset; // @[SynInMask.scala 83:42]
  wire  _T_174 = io_valid & _T_169; // @[SynInMask.scala 85:55]
  wire  _T_175 = _T_174 & noWait; // @[SynInMask.scala 85:92]
  wire  _T_177 = _T_175 & _T_162; // @[SynInMask.scala 85:102]
  wire  _T_178 = _T_177 & dmaCGRAInMask_1; // @[SynInMask.scala 85:122]
  reg [31:0] inDatasWire_1; // @[Reg.scala 27:20]
  wire  _T_182 = _T_169 & io_valid; // @[SynInMask.scala 86:90]
  wire  _T_183 = _T_182 & noWait; // @[SynInMask.scala 86:102]
  wire  _T_185 = _T_183 & _T_162; // @[SynInMask.scala 86:111]
  wire  _T_186 = _T_185 & dmaCGRAInMask_1; // @[SynInMask.scala 86:131]
  wire  _T_197 = ~_T_196; // @[SynInMask.scala 83:27]
  wire  _T_198 = dataRst & _T_197; // @[SynInMask.scala 83:24]
  wire  _T_200 = _T_198 | reset; // @[SynInMask.scala 83:42]
  wire  _T_207 = io_valid & _T_202; // @[SynInMask.scala 85:55]
  wire  _T_208 = _T_207 & noWait; // @[SynInMask.scala 85:92]
  wire  _T_210 = _T_208 & _T_195; // @[SynInMask.scala 85:102]
  wire  _T_211 = _T_210 & dmaCGRAInMask_2; // @[SynInMask.scala 85:122]
  reg [31:0] inDatasWire_2; // @[Reg.scala 27:20]
  wire  _T_215 = _T_202 & io_valid; // @[SynInMask.scala 86:90]
  wire  _T_216 = _T_215 & noWait; // @[SynInMask.scala 86:102]
  wire  _T_218 = _T_216 & _T_195; // @[SynInMask.scala 86:111]
  wire  _T_219 = _T_218 & dmaCGRAInMask_2; // @[SynInMask.scala 86:131]
  wire  _T_230 = ~_T_229; // @[SynInMask.scala 83:27]
  wire  _T_231 = dataRst & _T_230; // @[SynInMask.scala 83:24]
  wire  _T_233 = _T_231 | reset; // @[SynInMask.scala 83:42]
  wire  _T_240 = io_valid & _T_235; // @[SynInMask.scala 85:55]
  wire  _T_241 = _T_240 & noWait; // @[SynInMask.scala 85:92]
  wire  _T_243 = _T_241 & _T_228; // @[SynInMask.scala 85:102]
  wire  _T_244 = _T_243 & dmaCGRAInMask_3; // @[SynInMask.scala 85:122]
  reg [31:0] inDatasWire_3; // @[Reg.scala 27:20]
  wire  _T_248 = _T_235 & io_valid; // @[SynInMask.scala 86:90]
  wire  _T_249 = _T_248 & noWait; // @[SynInMask.scala 86:102]
  wire  _T_251 = _T_249 & _T_228; // @[SynInMask.scala 86:111]
  wire  _T_252 = _T_251 & dmaCGRAInMask_3; // @[SynInMask.scala 86:131]
  wire  _T_263 = ~_T_262; // @[SynInMask.scala 83:27]
  wire  _T_264 = dataRst & _T_263; // @[SynInMask.scala 83:24]
  wire  _T_266 = _T_264 | reset; // @[SynInMask.scala 83:42]
  wire  _T_273 = io_valid & _T_268; // @[SynInMask.scala 85:55]
  wire  _T_274 = _T_273 & noWait; // @[SynInMask.scala 85:92]
  wire  _T_276 = _T_274 & _T_261; // @[SynInMask.scala 85:102]
  wire  _T_277 = _T_276 & dmaCGRAInMask_4; // @[SynInMask.scala 85:122]
  reg [31:0] inDatasWire_4; // @[Reg.scala 27:20]
  wire  _T_281 = _T_268 & io_valid; // @[SynInMask.scala 86:90]
  wire  _T_282 = _T_281 & noWait; // @[SynInMask.scala 86:102]
  wire  _T_284 = _T_282 & _T_261; // @[SynInMask.scala 86:111]
  wire  _T_285 = _T_284 & dmaCGRAInMask_4; // @[SynInMask.scala 86:131]
  wire  _T_296 = ~_T_295; // @[SynInMask.scala 83:27]
  wire  _T_297 = dataRst & _T_296; // @[SynInMask.scala 83:24]
  wire  _T_299 = _T_297 | reset; // @[SynInMask.scala 83:42]
  wire  _T_306 = io_valid & _T_301; // @[SynInMask.scala 85:55]
  wire  _T_307 = _T_306 & noWait; // @[SynInMask.scala 85:92]
  wire  _T_309 = _T_307 & _T_294; // @[SynInMask.scala 85:102]
  wire  _T_310 = _T_309 & dmaCGRAInMask_5; // @[SynInMask.scala 85:122]
  reg [31:0] inDatasWire_5; // @[Reg.scala 27:20]
  wire  _T_314 = _T_301 & io_valid; // @[SynInMask.scala 86:90]
  wire  _T_315 = _T_314 & noWait; // @[SynInMask.scala 86:102]
  wire  _T_317 = _T_315 & _T_294; // @[SynInMask.scala 86:111]
  wire  _T_318 = _T_317 & dmaCGRAInMask_5; // @[SynInMask.scala 86:131]
  wire  _T_329 = ~_T_328; // @[SynInMask.scala 83:27]
  wire  _T_330 = dataRst & _T_329; // @[SynInMask.scala 83:24]
  wire  _T_332 = _T_330 | reset; // @[SynInMask.scala 83:42]
  wire  _T_339 = io_valid & _T_334; // @[SynInMask.scala 85:55]
  wire  _T_340 = _T_339 & noWait; // @[SynInMask.scala 85:92]
  wire  _T_342 = _T_340 & _T_327; // @[SynInMask.scala 85:102]
  wire  _T_343 = _T_342 & dmaCGRAInMask_6; // @[SynInMask.scala 85:122]
  reg [31:0] inDatasWire_6; // @[Reg.scala 27:20]
  wire  _T_347 = _T_334 & io_valid; // @[SynInMask.scala 86:90]
  wire  _T_348 = _T_347 & noWait; // @[SynInMask.scala 86:102]
  wire  _T_350 = _T_348 & _T_327; // @[SynInMask.scala 86:111]
  wire  _T_351 = _T_350 & dmaCGRAInMask_6; // @[SynInMask.scala 86:131]
  wire  _T_362 = ~_T_361; // @[SynInMask.scala 83:27]
  wire  _T_363 = dataRst & _T_362; // @[SynInMask.scala 83:24]
  wire  _T_365 = _T_363 | reset; // @[SynInMask.scala 83:42]
  wire  _T_372 = io_valid & _T_367; // @[SynInMask.scala 85:55]
  wire  _T_373 = _T_372 & noWait; // @[SynInMask.scala 85:92]
  wire  _T_375 = _T_373 & _T_360; // @[SynInMask.scala 85:102]
  wire  _T_376 = _T_375 & dmaCGRAInMask_7; // @[SynInMask.scala 85:122]
  reg [31:0] inDatasWire_7; // @[Reg.scala 27:20]
  wire  _T_380 = _T_367 & io_valid; // @[SynInMask.scala 86:90]
  wire  _T_381 = _T_380 & noWait; // @[SynInMask.scala 86:102]
  wire  _T_383 = _T_381 & _T_360; // @[SynInMask.scala 86:111]
  wire  _T_384 = _T_383 & dmaCGRAInMask_7; // @[SynInMask.scala 86:131]
  wire  _T_395 = ~_T_394; // @[SynInMask.scala 83:27]
  wire  _T_396 = dataRst & _T_395; // @[SynInMask.scala 83:24]
  wire  _T_398 = _T_396 | reset; // @[SynInMask.scala 83:42]
  wire  _T_405 = io_valid & _T_400; // @[SynInMask.scala 85:55]
  wire  _T_406 = _T_405 & noWait; // @[SynInMask.scala 85:92]
  wire  _T_408 = _T_406 & _T_393; // @[SynInMask.scala 85:102]
  wire  _T_409 = _T_408 & dmaCGRAInMask_8; // @[SynInMask.scala 85:122]
  reg [31:0] inDatasWire_8; // @[Reg.scala 27:20]
  wire  _T_413 = _T_400 & io_valid; // @[SynInMask.scala 86:90]
  wire  _T_414 = _T_413 & noWait; // @[SynInMask.scala 86:102]
  wire  _T_416 = _T_414 & _T_393; // @[SynInMask.scala 86:111]
  wire  _T_417 = _T_416 & dmaCGRAInMask_8; // @[SynInMask.scala 86:131]
  wire  _T_428 = ~_T_427; // @[SynInMask.scala 83:27]
  wire  _T_429 = dataRst & _T_428; // @[SynInMask.scala 83:24]
  wire  _T_431 = _T_429 | reset; // @[SynInMask.scala 83:42]
  wire  _T_438 = io_valid & _T_433; // @[SynInMask.scala 85:55]
  wire  _T_439 = _T_438 & noWait; // @[SynInMask.scala 85:92]
  wire  _T_441 = _T_439 & _T_426; // @[SynInMask.scala 85:102]
  wire  _T_442 = _T_441 & dmaCGRAInMask_9; // @[SynInMask.scala 85:122]
  reg [31:0] inDatasWire_9; // @[Reg.scala 27:20]
  wire  _T_446 = _T_433 & io_valid; // @[SynInMask.scala 86:90]
  wire  _T_447 = _T_446 & noWait; // @[SynInMask.scala 86:102]
  wire  _T_449 = _T_447 & _T_426; // @[SynInMask.scala 86:111]
  wire  _T_450 = _T_449 & dmaCGRAInMask_9; // @[SynInMask.scala 86:131]
  wire  _T_461 = ~_T_460; // @[SynInMask.scala 83:27]
  wire  _T_462 = dataRst & _T_461; // @[SynInMask.scala 83:24]
  wire  _T_464 = _T_462 | reset; // @[SynInMask.scala 83:42]
  wire  _T_471 = io_valid & _T_466; // @[SynInMask.scala 85:55]
  wire  _T_472 = _T_471 & noWait; // @[SynInMask.scala 85:92]
  wire  _T_474 = _T_472 & _T_459; // @[SynInMask.scala 85:102]
  wire  _T_475 = _T_474 & dmaCGRAInMask_10; // @[SynInMask.scala 85:122]
  reg [31:0] inDatasWire_10; // @[Reg.scala 27:20]
  wire  _T_479 = _T_466 & io_valid; // @[SynInMask.scala 86:90]
  wire  _T_480 = _T_479 & noWait; // @[SynInMask.scala 86:102]
  wire  _T_482 = _T_480 & _T_459; // @[SynInMask.scala 86:111]
  wire  _T_483 = _T_482 & dmaCGRAInMask_10; // @[SynInMask.scala 86:131]
  wire  _T_494 = ~_T_493; // @[SynInMask.scala 83:27]
  wire  _T_495 = dataRst & _T_494; // @[SynInMask.scala 83:24]
  wire  _T_497 = _T_495 | reset; // @[SynInMask.scala 83:42]
  wire  _T_504 = io_valid & _T_499; // @[SynInMask.scala 85:55]
  wire  _T_505 = _T_504 & noWait; // @[SynInMask.scala 85:92]
  wire  _T_507 = _T_505 & _T_492; // @[SynInMask.scala 85:102]
  wire  _T_508 = _T_507 & dmaCGRAInMask_11; // @[SynInMask.scala 85:122]
  reg [31:0] inDatasWire_11; // @[Reg.scala 27:20]
  wire  _T_512 = _T_499 & io_valid; // @[SynInMask.scala 86:90]
  wire  _T_513 = _T_512 & noWait; // @[SynInMask.scala 86:102]
  wire  _T_515 = _T_513 & _T_492; // @[SynInMask.scala 86:111]
  wire  _T_516 = _T_515 & dmaCGRAInMask_11; // @[SynInMask.scala 86:131]
  wire  _T_527 = ~_T_526; // @[SynInMask.scala 83:27]
  wire  _T_528 = dataRst & _T_527; // @[SynInMask.scala 83:24]
  wire  _T_530 = _T_528 | reset; // @[SynInMask.scala 83:42]
  wire  _T_537 = io_valid & _T_532; // @[SynInMask.scala 85:55]
  wire  _T_538 = _T_537 & noWait; // @[SynInMask.scala 85:92]
  wire  _T_540 = _T_538 & _T_525; // @[SynInMask.scala 85:102]
  wire  _T_541 = _T_540 & dmaCGRAInMask_12; // @[SynInMask.scala 85:122]
  reg [31:0] inDatasWire_12; // @[Reg.scala 27:20]
  wire  _T_545 = _T_532 & io_valid; // @[SynInMask.scala 86:90]
  wire  _T_546 = _T_545 & noWait; // @[SynInMask.scala 86:102]
  wire  _T_548 = _T_546 & _T_525; // @[SynInMask.scala 86:111]
  wire  _T_549 = _T_548 & dmaCGRAInMask_12; // @[SynInMask.scala 86:131]
  wire  _T_560 = ~_T_559; // @[SynInMask.scala 83:27]
  wire  _T_561 = dataRst & _T_560; // @[SynInMask.scala 83:24]
  wire  _T_563 = _T_561 | reset; // @[SynInMask.scala 83:42]
  wire  _T_570 = io_valid & _T_565; // @[SynInMask.scala 85:55]
  wire  _T_571 = _T_570 & noWait; // @[SynInMask.scala 85:92]
  wire  _T_573 = _T_571 & _T_558; // @[SynInMask.scala 85:102]
  wire  _T_574 = _T_573 & dmaCGRAInMask_13; // @[SynInMask.scala 85:122]
  reg [31:0] inDatasWire_13; // @[Reg.scala 27:20]
  wire  _T_578 = _T_565 & io_valid; // @[SynInMask.scala 86:90]
  wire  _T_579 = _T_578 & noWait; // @[SynInMask.scala 86:102]
  wire  _T_581 = _T_579 & _T_558; // @[SynInMask.scala 86:111]
  wire  _T_582 = _T_581 & dmaCGRAInMask_13; // @[SynInMask.scala 86:131]
  wire  _T_593 = ~_T_592; // @[SynInMask.scala 83:27]
  wire  _T_594 = dataRst & _T_593; // @[SynInMask.scala 83:24]
  wire  _T_596 = _T_594 | reset; // @[SynInMask.scala 83:42]
  wire  _T_603 = io_valid & _T_598; // @[SynInMask.scala 85:55]
  wire  _T_604 = _T_603 & noWait; // @[SynInMask.scala 85:92]
  wire  _T_606 = _T_604 & _T_591; // @[SynInMask.scala 85:102]
  wire  _T_607 = _T_606 & dmaCGRAInMask_14; // @[SynInMask.scala 85:122]
  reg [31:0] inDatasWire_14; // @[Reg.scala 27:20]
  wire  _T_611 = _T_598 & io_valid; // @[SynInMask.scala 86:90]
  wire  _T_612 = _T_611 & noWait; // @[SynInMask.scala 86:102]
  wire  _T_614 = _T_612 & _T_591; // @[SynInMask.scala 86:111]
  wire  _T_615 = _T_614 & dmaCGRAInMask_14; // @[SynInMask.scala 86:131]
  wire  _T_626 = ~_T_625; // @[SynInMask.scala 83:27]
  wire  _T_627 = dataRst & _T_626; // @[SynInMask.scala 83:24]
  wire  _T_629 = _T_627 | reset; // @[SynInMask.scala 83:42]
  wire  _T_636 = io_valid & _T_631; // @[SynInMask.scala 85:55]
  wire  _T_637 = _T_636 & noWait; // @[SynInMask.scala 85:92]
  wire  _T_639 = _T_637 & _T_624; // @[SynInMask.scala 85:102]
  wire  _T_640 = _T_639 & dmaCGRAInMask_15; // @[SynInMask.scala 85:122]
  reg [31:0] inDatasWire_15; // @[Reg.scala 27:20]
  wire  _T_644 = _T_631 & io_valid; // @[SynInMask.scala 86:90]
  wire  _T_645 = _T_644 & noWait; // @[SynInMask.scala 86:102]
  wire  _T_647 = _T_645 & _T_624; // @[SynInMask.scala 86:111]
  wire  _T_648 = _T_647 & dmaCGRAInMask_15; // @[SynInMask.scala 86:131]
  wire  _T_680 = dataRst & outValidsWire_0; // @[SynInMask.scala 105:33]
  wire  _T_681 = _T_680 & dmaEnWR_0; // @[SynInMask.scala 105:52]
  wire  _T_683 = dataRst & outValidsWire_1; // @[SynInMask.scala 105:33]
  wire  _T_684 = _T_683 & dmaEnWR_0; // @[SynInMask.scala 105:52]
  wire  _T_686 = dataRst & outValidsWire_2; // @[SynInMask.scala 105:33]
  wire  _T_687 = _T_686 & dmaEnWR_0; // @[SynInMask.scala 105:52]
  wire  _T_689 = dataRst & outValidsWire_3; // @[SynInMask.scala 105:33]
  wire  _T_690 = _T_689 & dmaEnWR_0; // @[SynInMask.scala 105:52]
  wire  _T_692 = dataRst & outValidsWire_4; // @[SynInMask.scala 105:33]
  wire  _T_693 = _T_692 & dmaEnWR_0; // @[SynInMask.scala 105:52]
  wire  _T_695 = dataRst & outValidsWire_5; // @[SynInMask.scala 105:33]
  wire  _T_696 = _T_695 & dmaEnWR_0; // @[SynInMask.scala 105:52]
  wire  _T_698 = dataRst & outValidsWire_6; // @[SynInMask.scala 105:33]
  wire  _T_699 = _T_698 & dmaEnWR_0; // @[SynInMask.scala 105:52]
  wire  _T_701 = dataRst & outValidsWire_7; // @[SynInMask.scala 105:33]
  wire  _T_702 = _T_701 & dmaEnWR_0; // @[SynInMask.scala 105:52]
  wire  _T_704 = dataRst & outValidsWire_8; // @[SynInMask.scala 105:33]
  wire  _T_705 = _T_704 & dmaEnWR_0; // @[SynInMask.scala 105:52]
  wire  _T_707 = dataRst & outValidsWire_9; // @[SynInMask.scala 105:33]
  wire  _T_708 = _T_707 & dmaEnWR_0; // @[SynInMask.scala 105:52]
  wire  _T_710 = dataRst & outValidsWire_10; // @[SynInMask.scala 105:33]
  wire  _T_711 = _T_710 & dmaEnWR_0; // @[SynInMask.scala 105:52]
  wire  _T_713 = dataRst & outValidsWire_11; // @[SynInMask.scala 105:33]
  wire  _T_714 = _T_713 & dmaEnWR_0; // @[SynInMask.scala 105:52]
  wire  _T_716 = dataRst & outValidsWire_12; // @[SynInMask.scala 105:33]
  wire  _T_717 = _T_716 & dmaEnWR_0; // @[SynInMask.scala 105:52]
  wire  _T_719 = dataRst & outValidsWire_13; // @[SynInMask.scala 105:33]
  wire  _T_720 = _T_719 & dmaEnWR_0; // @[SynInMask.scala 105:52]
  wire  _T_722 = dataRst & outValidsWire_14; // @[SynInMask.scala 105:33]
  wire  _T_723 = _T_722 & dmaEnWR_0; // @[SynInMask.scala 105:52]
  wire  _T_725 = dataRst & outValidsWire_15; // @[SynInMask.scala 105:33]
  wire  _T_726 = _T_725 & dmaEnWR_0; // @[SynInMask.scala 105:52]
  adressGenIn adrGenInst ( // @[SynInMask.scala 28:25]
    .clock(adrGenInst_clock),
    .reset(adrGenInst_reset),
    .io_validList_0(adrGenInst_io_validList_0),
    .io_validList_1(adrGenInst_io_validList_1),
    .io_validList_2(adrGenInst_io_validList_2),
    .io_validList_3(adrGenInst_io_validList_3),
    .io_validList_4(adrGenInst_io_validList_4),
    .io_validList_5(adrGenInst_io_validList_5),
    .io_validList_6(adrGenInst_io_validList_6),
    .io_validList_7(adrGenInst_io_validList_7),
    .io_validList_8(adrGenInst_io_validList_8),
    .io_validList_9(adrGenInst_io_validList_9),
    .io_validList_10(adrGenInst_io_validList_10),
    .io_validList_11(adrGenInst_io_validList_11),
    .io_validList_12(adrGenInst_io_validList_12),
    .io_validList_13(adrGenInst_io_validList_13),
    .io_validList_14(adrGenInst_io_validList_14),
    .io_update(adrGenInst_io_update),
    .io_clear(adrGenInst_io_clear),
    .io_sel1(adrGenInst_io_sel1),
    .io_sel2(adrGenInst_io_sel2)
  );
  assign io_ready = _T_678 ? readyList_15 : _T_677; // @[SynInMask.scala 97:12]
  assign io_dataOut_0 = {_T_681,inDatasWire_0}; // @[SynInMask.scala 105:19]
  assign io_dataOut_1 = {_T_684,inDatasWire_1}; // @[SynInMask.scala 105:19]
  assign io_dataOut_2 = {_T_687,inDatasWire_2}; // @[SynInMask.scala 105:19]
  assign io_dataOut_3 = {_T_690,inDatasWire_3}; // @[SynInMask.scala 105:19]
  assign io_dataOut_4 = {_T_693,inDatasWire_4}; // @[SynInMask.scala 105:19]
  assign io_dataOut_5 = {_T_696,inDatasWire_5}; // @[SynInMask.scala 105:19]
  assign io_dataOut_6 = {_T_699,inDatasWire_6}; // @[SynInMask.scala 105:19]
  assign io_dataOut_7 = {_T_702,inDatasWire_7}; // @[SynInMask.scala 105:19]
  assign io_dataOut_8 = {_T_705,inDatasWire_8}; // @[SynInMask.scala 105:19]
  assign io_dataOut_9 = {_T_708,inDatasWire_9}; // @[SynInMask.scala 105:19]
  assign io_dataOut_10 = {_T_711,inDatasWire_10}; // @[SynInMask.scala 105:19]
  assign io_dataOut_11 = {_T_714,inDatasWire_11}; // @[SynInMask.scala 105:19]
  assign io_dataOut_12 = {_T_717,inDatasWire_12}; // @[SynInMask.scala 105:19]
  assign io_dataOut_13 = {_T_720,inDatasWire_13}; // @[SynInMask.scala 105:19]
  assign io_dataOut_14 = {_T_723,inDatasWire_14}; // @[SynInMask.scala 105:19]
  assign io_dataOut_15 = {_T_726,inDatasWire_15}; // @[SynInMask.scala 105:19]
  assign adrGenInst_clock = clock;
  assign adrGenInst_reset = reset;
  assign adrGenInst_io_validList_0 = dmaCtrl_0[64]; // @[SynInMask.scala 51:27]
  assign adrGenInst_io_validList_1 = dmaCtrl_0[65]; // @[SynInMask.scala 51:27]
  assign adrGenInst_io_validList_2 = dmaCtrl_0[66]; // @[SynInMask.scala 51:27]
  assign adrGenInst_io_validList_3 = dmaCtrl_0[67]; // @[SynInMask.scala 51:27]
  assign adrGenInst_io_validList_4 = dmaCtrl_0[68]; // @[SynInMask.scala 51:27]
  assign adrGenInst_io_validList_5 = dmaCtrl_0[69]; // @[SynInMask.scala 51:27]
  assign adrGenInst_io_validList_6 = dmaCtrl_0[70]; // @[SynInMask.scala 51:27]
  assign adrGenInst_io_validList_7 = dmaCtrl_0[71]; // @[SynInMask.scala 51:27]
  assign adrGenInst_io_validList_8 = dmaCtrl_0[72]; // @[SynInMask.scala 51:27]
  assign adrGenInst_io_validList_9 = dmaCtrl_0[73]; // @[SynInMask.scala 51:27]
  assign adrGenInst_io_validList_10 = dmaCtrl_0[74]; // @[SynInMask.scala 51:27]
  assign adrGenInst_io_validList_11 = dmaCtrl_0[75]; // @[SynInMask.scala 51:27]
  assign adrGenInst_io_validList_12 = dmaCtrl_0[76]; // @[SynInMask.scala 51:27]
  assign adrGenInst_io_validList_13 = dmaCtrl_0[77]; // @[SynInMask.scala 51:27]
  assign adrGenInst_io_validList_14 = dmaCtrl_0[78]; // @[SynInMask.scala 51:27]
  assign adrGenInst_io_update = readySel & io_valid; // @[SynInMask.scala 49:24]
  assign adrGenInst_io_clear = clearUp & updateWire; // @[SynInMask.scala 50:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  clearCountReg = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  outValidsWire_15 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  outValidsWire_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  outValidsWire_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  outValidsWire_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  outValidsWire_3 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  outValidsWire_4 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  outValidsWire_5 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  outValidsWire_6 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  outValidsWire_7 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  outValidsWire_8 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  outValidsWire_9 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  outValidsWire_10 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  outValidsWire_11 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  outValidsWire_12 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  outValidsWire_13 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  outValidsWire_14 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  delayCnt = _RAND_17[5:0];
  _RAND_18 = {1{`RANDOM}};
  delayReg = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  inDatasWire_0 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  inDatasWire_1 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  inDatasWire_2 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  inDatasWire_3 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  inDatasWire_4 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  inDatasWire_5 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  inDatasWire_6 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  inDatasWire_7 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  inDatasWire_8 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  inDatasWire_9 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  inDatasWire_10 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  inDatasWire_11 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  inDatasWire_12 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  inDatasWire_13 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  inDatasWire_14 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  inDatasWire_15 = _RAND_34[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      clearCountReg <= 4'h0;
    end else if (updateWire) begin
      if (clearUp) begin
        clearCountReg <= 4'h0;
      end else begin
        clearCountReg <= _T_71;
      end
    end
    if (_T_629) begin
      outValidsWire_15 <= 1'h0;
    end else if (_T_648) begin
      outValidsWire_15 <= io_valid;
    end
    if (_T_134) begin
      outValidsWire_0 <= 1'h0;
    end else if (_T_153) begin
      outValidsWire_0 <= io_valid;
    end
    if (_T_167) begin
      outValidsWire_1 <= 1'h0;
    end else if (_T_186) begin
      outValidsWire_1 <= io_valid;
    end
    if (_T_200) begin
      outValidsWire_2 <= 1'h0;
    end else if (_T_219) begin
      outValidsWire_2 <= io_valid;
    end
    if (_T_233) begin
      outValidsWire_3 <= 1'h0;
    end else if (_T_252) begin
      outValidsWire_3 <= io_valid;
    end
    if (_T_266) begin
      outValidsWire_4 <= 1'h0;
    end else if (_T_285) begin
      outValidsWire_4 <= io_valid;
    end
    if (_T_299) begin
      outValidsWire_5 <= 1'h0;
    end else if (_T_318) begin
      outValidsWire_5 <= io_valid;
    end
    if (_T_332) begin
      outValidsWire_6 <= 1'h0;
    end else if (_T_351) begin
      outValidsWire_6 <= io_valid;
    end
    if (_T_365) begin
      outValidsWire_7 <= 1'h0;
    end else if (_T_384) begin
      outValidsWire_7 <= io_valid;
    end
    if (_T_398) begin
      outValidsWire_8 <= 1'h0;
    end else if (_T_417) begin
      outValidsWire_8 <= io_valid;
    end
    if (_T_431) begin
      outValidsWire_9 <= 1'h0;
    end else if (_T_450) begin
      outValidsWire_9 <= io_valid;
    end
    if (_T_464) begin
      outValidsWire_10 <= 1'h0;
    end else if (_T_483) begin
      outValidsWire_10 <= io_valid;
    end
    if (_T_497) begin
      outValidsWire_11 <= 1'h0;
    end else if (_T_516) begin
      outValidsWire_11 <= io_valid;
    end
    if (_T_530) begin
      outValidsWire_12 <= 1'h0;
    end else if (_T_549) begin
      outValidsWire_12 <= io_valid;
    end
    if (_T_563) begin
      outValidsWire_13 <= 1'h0;
    end else if (_T_582) begin
      outValidsWire_13 <= io_valid;
    end
    if (_T_596) begin
      outValidsWire_14 <= 1'h0;
    end else if (_T_615) begin
      outValidsWire_14 <= io_valid;
    end
    if (reset) begin
      delayCnt <= 6'h0;
    end else if (_T_120) begin
      if (_T_116) begin
        delayCnt <= _T_118;
      end else begin
        delayCnt <= 6'h0;
      end
    end
    if (reset) begin
      delayReg <= 6'h0;
    end else if (io_delayen) begin
      delayReg <= io_delayCycle[5:0];
    end
    if (_T_134) begin
      inDatasWire_0 <= 32'h0;
    end else if (_T_145) begin
      if (_T_122) begin
        inDatasWire_0 <= io_dataIn[31:0];
      end else begin
        inDatasWire_0 <= io_dataIn[63:32];
      end
    end
    if (_T_167) begin
      inDatasWire_1 <= 32'h0;
    end else if (_T_178) begin
      if (_T_650) begin
        inDatasWire_1 <= io_dataIn[31:0];
      end else begin
        inDatasWire_1 <= io_dataIn[63:32];
      end
    end
    if (_T_200) begin
      inDatasWire_2 <= 32'h0;
    end else if (_T_211) begin
      if (_T_652) begin
        inDatasWire_2 <= io_dataIn[31:0];
      end else begin
        inDatasWire_2 <= io_dataIn[63:32];
      end
    end
    if (_T_233) begin
      inDatasWire_3 <= 32'h0;
    end else if (_T_244) begin
      if (_T_654) begin
        inDatasWire_3 <= io_dataIn[31:0];
      end else begin
        inDatasWire_3 <= io_dataIn[63:32];
      end
    end
    if (_T_266) begin
      inDatasWire_4 <= 32'h0;
    end else if (_T_277) begin
      if (_T_656) begin
        inDatasWire_4 <= io_dataIn[31:0];
      end else begin
        inDatasWire_4 <= io_dataIn[63:32];
      end
    end
    if (_T_299) begin
      inDatasWire_5 <= 32'h0;
    end else if (_T_310) begin
      if (_T_658) begin
        inDatasWire_5 <= io_dataIn[31:0];
      end else begin
        inDatasWire_5 <= io_dataIn[63:32];
      end
    end
    if (_T_332) begin
      inDatasWire_6 <= 32'h0;
    end else if (_T_343) begin
      if (_T_660) begin
        inDatasWire_6 <= io_dataIn[31:0];
      end else begin
        inDatasWire_6 <= io_dataIn[63:32];
      end
    end
    if (_T_365) begin
      inDatasWire_7 <= 32'h0;
    end else if (_T_376) begin
      if (_T_662) begin
        inDatasWire_7 <= io_dataIn[31:0];
      end else begin
        inDatasWire_7 <= io_dataIn[63:32];
      end
    end
    if (_T_398) begin
      inDatasWire_8 <= 32'h0;
    end else if (_T_409) begin
      if (_T_664) begin
        inDatasWire_8 <= io_dataIn[31:0];
      end else begin
        inDatasWire_8 <= io_dataIn[63:32];
      end
    end
    if (_T_431) begin
      inDatasWire_9 <= 32'h0;
    end else if (_T_442) begin
      if (_T_666) begin
        inDatasWire_9 <= io_dataIn[31:0];
      end else begin
        inDatasWire_9 <= io_dataIn[63:32];
      end
    end
    if (_T_464) begin
      inDatasWire_10 <= 32'h0;
    end else if (_T_475) begin
      if (_T_668) begin
        inDatasWire_10 <= io_dataIn[31:0];
      end else begin
        inDatasWire_10 <= io_dataIn[63:32];
      end
    end
    if (_T_497) begin
      inDatasWire_11 <= 32'h0;
    end else if (_T_508) begin
      if (_T_670) begin
        inDatasWire_11 <= io_dataIn[31:0];
      end else begin
        inDatasWire_11 <= io_dataIn[63:32];
      end
    end
    if (_T_530) begin
      inDatasWire_12 <= 32'h0;
    end else if (_T_541) begin
      if (_T_672) begin
        inDatasWire_12 <= io_dataIn[31:0];
      end else begin
        inDatasWire_12 <= io_dataIn[63:32];
      end
    end
    if (_T_563) begin
      inDatasWire_13 <= 32'h0;
    end else if (_T_574) begin
      if (_T_674) begin
        inDatasWire_13 <= io_dataIn[31:0];
      end else begin
        inDatasWire_13 <= io_dataIn[63:32];
      end
    end
    if (_T_596) begin
      inDatasWire_14 <= 32'h0;
    end else if (_T_607) begin
      if (_T_676) begin
        inDatasWire_14 <= io_dataIn[31:0];
      end else begin
        inDatasWire_14 <= io_dataIn[63:32];
      end
    end
    if (_T_629) begin
      inDatasWire_15 <= 32'h0;
    end else if (_T_640) begin
      if (_T_678) begin
        inDatasWire_15 <= io_dataIn[31:0];
      end else begin
        inDatasWire_15 <= io_dataIn[63:32];
      end
    end
  end
endmodule
module Mul(
  input         clock,
  input         reset,
  input         io_mulValid,
  input  [31:0] io_multiplicand,
  input  [31:0] io_multiplier,
  output        io_outValid,
  output [31:0] io_resultLow
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  _T; // @[Mul.scala 40:26]
  wire [63:0] _T_1 = io_multiplicand * io_multiplier; // @[Mul.scala 41:39]
  reg [63:0] _T_2; // @[Mul.scala 41:22]
  assign io_outValid = _T; // @[Mul.scala 40:17]
  assign io_resultLow = _T_2[31:0]; // @[Mul.scala 42:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  _T_2 = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T <= 1'h0;
    end else begin
      _T <= io_mulValid;
    end
    if (reset) begin
      _T_2 <= 64'h0;
    end else begin
      _T_2 <= _T_1;
    end
  end
endmodule
module Acc(
  input         clock,
  input         reset,
  input  [7:0]  io_iniVal,
  input  [7:0]  io_counter,
  input  [32:0] io_inputVal,
  output [32:0] io_outputVal
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  valid = io_inputVal[32]; // @[Acc.scala 12:26]
  wire [31:0] inVal = io_inputVal[31:0]; // @[Acc.scala 13:26]
  reg [7:0] accCntReg; // @[Reg.scala 27:20]
  wire  cntFinish = accCntReg == io_counter; // @[Acc.scala 15:30]
  wire [7:0] _T_3 = accCntReg + 8'h1; // @[Acc.scala 24:18]
  wire  _T_5 = valid | cntFinish; // @[Acc.scala 26:16]
  wire  _T_6 = accCntReg == 8'h0; // @[Acc.scala 34:31]
  wire  _T_7 = cntFinish | _T_6; // @[Acc.scala 34:18]
  wire [31:0] _GEN_2 = {{24'd0}, io_iniVal}; // @[Acc.scala 35:15]
  wire [31:0] _T_9 = inVal + _GEN_2; // @[Acc.scala 35:15]
  reg [31:0] accValReg; // @[Reg.scala 27:20]
  wire [31:0] _T_11 = inVal + accValReg; // @[Acc.scala 36:15]
  wire [31:0] _T_15 = cntFinish ? accValReg : 32'h0; // @[Acc.scala 49:8]
  assign io_outputVal = {cntFinish,_T_15}; // @[Acc.scala 47:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  accCntReg = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  accValReg = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      accCntReg <= 8'h0;
    end else if (_T_5) begin
      if (cntFinish) begin
        accCntReg <= {{7'd0}, valid};
      end else begin
        accCntReg <= _T_3;
      end
    end
    if (reset) begin
      accValReg <= 32'h0;
    end else if (_T_5) begin
      if (valid) begin
        if (_T_7) begin
          accValReg <= _T_9;
        end else begin
          accValReg <= _T_11;
        end
      end else begin
        accValReg <= 32'h0;
      end
    end
  end
endmodule
module ALU0(
  input         clock,
  input         reset,
  input  [20:0] io_cfg,
  input  [32:0] io_inputs_0,
  input  [32:0] io_inputs_1,
  output [32:0] io_outputs_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  Mul_clock; // @[ALU.scala 88:30]
  wire  Mul_reset; // @[ALU.scala 88:30]
  wire  Mul_io_mulValid; // @[ALU.scala 88:30]
  wire [31:0] Mul_io_multiplicand; // @[ALU.scala 88:30]
  wire [31:0] Mul_io_multiplier; // @[ALU.scala 88:30]
  wire  Mul_io_outValid; // @[ALU.scala 88:30]
  wire [31:0] Mul_io_resultLow; // @[ALU.scala 88:30]
  wire  Acc_clock; // @[ALU.scala 116:32]
  wire  Acc_reset; // @[ALU.scala 116:32]
  wire [7:0] Acc_io_iniVal; // @[ALU.scala 116:32]
  wire [7:0] Acc_io_counter; // @[ALU.scala 116:32]
  wire [32:0] Acc_io_inputVal; // @[ALU.scala 116:32]
  wire [32:0] Acc_io_outputVal; // @[ALU.scala 116:32]
  reg [32:0] inputsWire_0; // @[Reg.scala 27:20]
  reg [32:0] inputsWire_1; // @[Reg.scala 27:20]
  wire  _T_2 = inputsWire_0[32] & inputsWire_1[32]; // @[ALU.scala 39:41]
  wire  _T_17 = 5'h1 == io_cfg[4:0]; // @[Mux.scala 80:60]
  wire  _T_18 = _T_17 & _T_2; // @[Mux.scala 80:57]
  wire  _T_19 = 5'h2 == io_cfg[4:0]; // @[Mux.scala 80:60]
  wire  _T_20 = _T_19 ? _T_2 : _T_18; // @[Mux.scala 80:57]
  wire  _T_21 = 5'h3 == io_cfg[4:0]; // @[Mux.scala 80:60]
  wire  _T_22 = _T_21 ? _T_2 : _T_20; // @[Mux.scala 80:57]
  wire  _T_23 = 5'h6 == io_cfg[4:0]; // @[Mux.scala 80:60]
  wire  _T_24 = _T_23 ? _T_2 : _T_22; // @[Mux.scala 80:57]
  wire  _T_25 = 5'h7 == io_cfg[4:0]; // @[Mux.scala 80:60]
  wire  _T_26 = _T_25 ? _T_2 : _T_24; // @[Mux.scala 80:57]
  wire  _T_27 = 5'h10 == io_cfg[4:0]; // @[Mux.scala 80:60]
  wire  en = _T_27 ? inputsWire_0[32] : _T_26; // @[Mux.scala 80:57]
  wire  _T_29 = ~io_inputs_0[32]; // @[ALU.scala 71:25]
  wire  _T_30 = en & _T_29; // @[ALU.scala 71:22]
  wire  _T_32 = _T_30 | reset; // @[ALU.scala 71:47]
  wire  _T_36 = ~io_inputs_1[32]; // @[ALU.scala 71:25]
  wire  _T_37 = en & _T_36; // @[ALU.scala 71:22]
  wire  _T_39 = _T_37 | reset; // @[ALU.scala 71:47]
  wire [31:0] _T_45 = inputsWire_0[31:0] + inputsWire_1[31:0]; // @[ALU.scala 85:62]
  wire [32:0] _T_46 = {en,_T_45}; // @[Cat.scala 29:58]
  wire [31:0] _T_50 = inputsWire_0[31:0] - inputsWire_1[31:0]; // @[ALU.scala 86:62]
  wire [32:0] _T_51 = {en,_T_50}; // @[Cat.scala 29:58]
  wire  _T_53 = io_cfg[4:0] == 5'h3; // @[ALU.scala 89:76]
  wire [32:0] _T_57 = {Mul_io_outValid,Mul_io_resultLow}; // @[Cat.scala 29:58]
  wire [31:0] _T_60 = inputsWire_0[31:0] | inputsWire_1[31:0]; // @[ALU.scala 104:61]
  wire [32:0] _T_61 = {en,_T_60}; // @[Cat.scala 29:58]
  wire [31:0] _T_64 = inputsWire_0[31:0] ^ inputsWire_1[31:0]; // @[ALU.scala 105:62]
  wire [32:0] _T_65 = {en,_T_64}; // @[Cat.scala 29:58]
  reg [32:0] _T_68; // @[ALU.scala 119:41]
  wire [32:0] _T_71 = _T_17 ? _T_46 : 33'h0; // @[Mux.scala 80:57]
  wire [32:0] _T_73 = _T_19 ? _T_51 : _T_71; // @[Mux.scala 80:57]
  wire [32:0] _T_75 = _T_21 ? _T_57 : _T_73; // @[Mux.scala 80:57]
  wire [32:0] _T_77 = _T_23 ? _T_61 : _T_75; // @[Mux.scala 80:57]
  wire [32:0] _T_79 = _T_25 ? _T_65 : _T_77; // @[Mux.scala 80:57]
  Mul Mul ( // @[ALU.scala 88:30]
    .clock(Mul_clock),
    .reset(Mul_reset),
    .io_mulValid(Mul_io_mulValid),
    .io_multiplicand(Mul_io_multiplicand),
    .io_multiplier(Mul_io_multiplier),
    .io_outValid(Mul_io_outValid),
    .io_resultLow(Mul_io_resultLow)
  );
  Acc Acc ( // @[ALU.scala 116:32]
    .clock(Acc_clock),
    .reset(Acc_reset),
    .io_iniVal(Acc_io_iniVal),
    .io_counter(Acc_io_counter),
    .io_inputVal(Acc_io_inputVal),
    .io_outputVal(Acc_io_outputVal)
  );
  assign io_outputs_0 = _T_27 ? Acc_io_outputVal : _T_79; // @[ALU.scala 129:16]
  assign Mul_clock = clock;
  assign Mul_reset = reset;
  assign Mul_io_mulValid = en & _T_53; // @[ALU.scala 89:30]
  assign Mul_io_multiplicand = inputsWire_0[31:0]; // @[ALU.scala 91:34]
  assign Mul_io_multiplier = inputsWire_1[31:0]; // @[ALU.scala 92:32]
  assign Acc_clock = clock;
  assign Acc_reset = reset;
  assign Acc_io_iniVal = io_cfg[20:13]; // @[ALU.scala 118:30]
  assign Acc_io_counter = io_cfg[12:5]; // @[ALU.scala 117:31]
  assign Acc_io_inputVal = _T_68; // @[ALU.scala 119:32]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  inputsWire_0 = _RAND_0[32:0];
  _RAND_1 = {2{`RANDOM}};
  inputsWire_1 = _RAND_1[32:0];
  _RAND_2 = {2{`RANDOM}};
  _T_68 = _RAND_2[32:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_32) begin
      inputsWire_0 <= 33'h0;
    end else if (io_inputs_0[32]) begin
      inputsWire_0 <= io_inputs_0;
    end
    if (_T_39) begin
      inputsWire_1 <= 33'h0;
    end else if (io_inputs_1[32]) begin
      inputsWire_1 <= io_inputs_1;
    end
    if (reset) begin
      _T_68 <= 33'h0;
    end else begin
      _T_68 <= io_inputs_0;
    end
  end
endmodule
module CfgMem(
  input         clock,
  input         reset,
  input         io_cfgEn,
  input  [31:0] io_cfgData,
  output [20:0] io_cfgOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] outWire_0; // @[Reg.scala 27:20]
  assign io_cfgOut = outWire_0[20:0]; // @[CfgMem.scala 22:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  outWire_0 = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      outWire_0 <= 32'h0;
    end else if (io_cfgEn) begin
      outWire_0 <= io_cfgData;
    end
  end
endmodule
module PE0(
  input         clock,
  input         reset,
  input         io_cfgEn,
  input  [31:0] io_cfgData,
  input  [32:0] io_inputs_0,
  input  [32:0] io_inputs_1,
  output [32:0] io_outputs_0
);
  wire  ALU0_clock; // @[TopModule.scala 186:48]
  wire  ALU0_reset; // @[TopModule.scala 186:48]
  wire [20:0] ALU0_io_cfg; // @[TopModule.scala 186:48]
  wire [32:0] ALU0_io_inputs_0; // @[TopModule.scala 186:48]
  wire [32:0] ALU0_io_inputs_1; // @[TopModule.scala 186:48]
  wire [32:0] ALU0_io_outputs_0; // @[TopModule.scala 186:48]
  wire  CfgMem_clock; // @[TopModule.scala 232:29]
  wire  CfgMem_reset; // @[TopModule.scala 232:29]
  wire  CfgMem_io_cfgEn; // @[TopModule.scala 232:29]
  wire [31:0] CfgMem_io_cfgData; // @[TopModule.scala 232:29]
  wire [20:0] CfgMem_io_cfgOut; // @[TopModule.scala 232:29]
  ALU0 ALU0 ( // @[TopModule.scala 186:48]
    .clock(ALU0_clock),
    .reset(ALU0_reset),
    .io_cfg(ALU0_io_cfg),
    .io_inputs_0(ALU0_io_inputs_0),
    .io_inputs_1(ALU0_io_inputs_1),
    .io_outputs_0(ALU0_io_outputs_0)
  );
  CfgMem CfgMem ( // @[TopModule.scala 232:29]
    .clock(CfgMem_clock),
    .reset(CfgMem_reset),
    .io_cfgEn(CfgMem_io_cfgEn),
    .io_cfgData(CfgMem_io_cfgData),
    .io_cfgOut(CfgMem_io_cfgOut)
  );
  assign io_outputs_0 = ALU0_io_outputs_0; // @[TopModule.scala 392:22]
  assign ALU0_clock = clock;
  assign ALU0_reset = reset;
  assign ALU0_io_cfg = CfgMem_io_cfgOut; // @[TopModule.scala 258:82]
  assign ALU0_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign ALU0_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign CfgMem_clock = clock;
  assign CfgMem_reset = reset;
  assign CfgMem_io_cfgEn = io_cfgEn; // @[TopModule.scala 239:34]
  assign CfgMem_io_cfgData = io_cfgData; // @[TopModule.scala 248:28]
endmodule
module ConstUnit0(
  input  [31:0] io_cfg,
  output [32:0] io_outputs_0
);
  assign io_outputs_0 = {1'h1,io_cfg}; // @[ConstUnit.scala 14:17]
endmodule
module MUX0(
  input  [4:0]  io_cfg,
  input  [32:0] io_inputs_0,
  input  [32:0] io_inputs_1,
  input  [32:0] io_inputs_2,
  input  [32:0] io_inputs_3,
  input  [32:0] io_inputs_4,
  input  [32:0] io_inputs_5,
  input  [32:0] io_inputs_6,
  input  [32:0] io_inputs_7,
  input  [32:0] io_inputs_8,
  input  [32:0] io_inputs_9,
  input  [32:0] io_inputs_10,
  input  [32:0] io_inputs_11,
  input  [32:0] io_inputs_12,
  input  [32:0] io_inputs_13,
  input  [32:0] io_inputs_14,
  input  [32:0] io_inputs_15,
  input  [32:0] io_inputs_16,
  output [32:0] io_outputs_0
);
  wire  _T = 5'h0 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_1 = _T ? io_inputs_0 : 33'h0; // @[Mux.scala 80:57]
  wire  _T_2 = 5'h1 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_3 = _T_2 ? io_inputs_1 : _T_1; // @[Mux.scala 80:57]
  wire  _T_4 = 5'h2 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_5 = _T_4 ? io_inputs_2 : _T_3; // @[Mux.scala 80:57]
  wire  _T_6 = 5'h3 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_7 = _T_6 ? io_inputs_3 : _T_5; // @[Mux.scala 80:57]
  wire  _T_8 = 5'h4 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_9 = _T_8 ? io_inputs_4 : _T_7; // @[Mux.scala 80:57]
  wire  _T_10 = 5'h5 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_11 = _T_10 ? io_inputs_5 : _T_9; // @[Mux.scala 80:57]
  wire  _T_12 = 5'h6 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_13 = _T_12 ? io_inputs_6 : _T_11; // @[Mux.scala 80:57]
  wire  _T_14 = 5'h7 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_15 = _T_14 ? io_inputs_7 : _T_13; // @[Mux.scala 80:57]
  wire  _T_16 = 5'h8 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_17 = _T_16 ? io_inputs_8 : _T_15; // @[Mux.scala 80:57]
  wire  _T_18 = 5'h9 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_19 = _T_18 ? io_inputs_9 : _T_17; // @[Mux.scala 80:57]
  wire  _T_20 = 5'ha == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_21 = _T_20 ? io_inputs_10 : _T_19; // @[Mux.scala 80:57]
  wire  _T_22 = 5'hb == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_23 = _T_22 ? io_inputs_11 : _T_21; // @[Mux.scala 80:57]
  wire  _T_24 = 5'hc == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_25 = _T_24 ? io_inputs_12 : _T_23; // @[Mux.scala 80:57]
  wire  _T_26 = 5'hd == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_27 = _T_26 ? io_inputs_13 : _T_25; // @[Mux.scala 80:57]
  wire  _T_28 = 5'he == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_29 = _T_28 ? io_inputs_14 : _T_27; // @[Mux.scala 80:57]
  wire  _T_30 = 5'hf == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_31 = _T_30 ? io_inputs_15 : _T_29; // @[Mux.scala 80:57]
  wire  _T_32 = 5'h10 == io_cfg; // @[Mux.scala 80:60]
  assign io_outputs_0 = _T_32 ? io_inputs_16 : _T_31; // @[Multiplexer.scala 16:17]
endmodule
module MUX8(
  input  [4:0]  io_cfg,
  input  [32:0] io_inputs_0,
  input  [32:0] io_inputs_1,
  input  [32:0] io_inputs_2,
  input  [32:0] io_inputs_3,
  input  [32:0] io_inputs_4,
  input  [32:0] io_inputs_5,
  input  [32:0] io_inputs_6,
  input  [32:0] io_inputs_7,
  input  [32:0] io_inputs_8,
  input  [32:0] io_inputs_9,
  input  [32:0] io_inputs_10,
  input  [32:0] io_inputs_11,
  input  [32:0] io_inputs_12,
  input  [32:0] io_inputs_13,
  input  [32:0] io_inputs_14,
  input  [32:0] io_inputs_15,
  input  [32:0] io_inputs_16,
  input  [32:0] io_inputs_17,
  output [32:0] io_outputs_0
);
  wire  _T = 5'h0 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_1 = _T ? io_inputs_0 : 33'h0; // @[Mux.scala 80:57]
  wire  _T_2 = 5'h1 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_3 = _T_2 ? io_inputs_1 : _T_1; // @[Mux.scala 80:57]
  wire  _T_4 = 5'h2 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_5 = _T_4 ? io_inputs_2 : _T_3; // @[Mux.scala 80:57]
  wire  _T_6 = 5'h3 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_7 = _T_6 ? io_inputs_3 : _T_5; // @[Mux.scala 80:57]
  wire  _T_8 = 5'h4 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_9 = _T_8 ? io_inputs_4 : _T_7; // @[Mux.scala 80:57]
  wire  _T_10 = 5'h5 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_11 = _T_10 ? io_inputs_5 : _T_9; // @[Mux.scala 80:57]
  wire  _T_12 = 5'h6 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_13 = _T_12 ? io_inputs_6 : _T_11; // @[Mux.scala 80:57]
  wire  _T_14 = 5'h7 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_15 = _T_14 ? io_inputs_7 : _T_13; // @[Mux.scala 80:57]
  wire  _T_16 = 5'h8 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_17 = _T_16 ? io_inputs_8 : _T_15; // @[Mux.scala 80:57]
  wire  _T_18 = 5'h9 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_19 = _T_18 ? io_inputs_9 : _T_17; // @[Mux.scala 80:57]
  wire  _T_20 = 5'ha == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_21 = _T_20 ? io_inputs_10 : _T_19; // @[Mux.scala 80:57]
  wire  _T_22 = 5'hb == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_23 = _T_22 ? io_inputs_11 : _T_21; // @[Mux.scala 80:57]
  wire  _T_24 = 5'hc == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_25 = _T_24 ? io_inputs_12 : _T_23; // @[Mux.scala 80:57]
  wire  _T_26 = 5'hd == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_27 = _T_26 ? io_inputs_13 : _T_25; // @[Mux.scala 80:57]
  wire  _T_28 = 5'he == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_29 = _T_28 ? io_inputs_14 : _T_27; // @[Mux.scala 80:57]
  wire  _T_30 = 5'hf == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_31 = _T_30 ? io_inputs_15 : _T_29; // @[Mux.scala 80:57]
  wire  _T_32 = 5'h10 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_33 = _T_32 ? io_inputs_16 : _T_31; // @[Mux.scala 80:57]
  wire  _T_34 = 5'h11 == io_cfg; // @[Mux.scala 80:60]
  assign io_outputs_0 = _T_34 ? io_inputs_17 : _T_33; // @[Multiplexer.scala 16:17]
endmodule
module MUXR0(
  input         clock,
  input         reset,
  input  [4:0]  io_cfg,
  input  [32:0] io_inputs_0,
  input  [32:0] io_inputs_1,
  input  [32:0] io_inputs_2,
  input  [32:0] io_inputs_3,
  input  [32:0] io_inputs_4,
  input  [32:0] io_inputs_5,
  input  [32:0] io_inputs_6,
  input  [32:0] io_inputs_7,
  input  [32:0] io_inputs_8,
  input  [32:0] io_inputs_9,
  input  [32:0] io_inputs_10,
  input  [32:0] io_inputs_11,
  input  [32:0] io_inputs_12,
  input  [32:0] io_inputs_13,
  input  [32:0] io_inputs_14,
  input  [32:0] io_inputs_15,
  input  [32:0] io_inputs_16,
  output [32:0] io_outputs_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _T = 5'h0 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_2 = 5'h1 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_4 = 5'h2 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_6 = 5'h3 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_8 = 5'h4 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_10 = 5'h5 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_12 = 5'h6 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_14 = 5'h7 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_16 = 5'h8 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_18 = 5'h9 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_20 = 5'ha == io_cfg; // @[Mux.scala 80:60]
  wire  _T_22 = 5'hb == io_cfg; // @[Mux.scala 80:60]
  wire  _T_24 = 5'hc == io_cfg; // @[Mux.scala 80:60]
  wire  _T_26 = 5'hd == io_cfg; // @[Mux.scala 80:60]
  wire  _T_28 = 5'he == io_cfg; // @[Mux.scala 80:60]
  wire  _T_30 = 5'hf == io_cfg; // @[Mux.scala 80:60]
  wire  _T_32 = 5'h10 == io_cfg; // @[Mux.scala 80:60]
  reg [32:0] _T_34; // @[MultiplexerR.scala 16:27]
  assign io_outputs_0 = _T_34; // @[MultiplexerR.scala 16:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_34 = _RAND_0[32:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_34 <= 33'h0;
    end else if (_T_32) begin
      _T_34 <= io_inputs_16;
    end else if (_T_30) begin
      _T_34 <= io_inputs_15;
    end else if (_T_28) begin
      _T_34 <= io_inputs_14;
    end else if (_T_26) begin
      _T_34 <= io_inputs_13;
    end else if (_T_24) begin
      _T_34 <= io_inputs_12;
    end else if (_T_22) begin
      _T_34 <= io_inputs_11;
    end else if (_T_20) begin
      _T_34 <= io_inputs_10;
    end else if (_T_18) begin
      _T_34 <= io_inputs_9;
    end else if (_T_16) begin
      _T_34 <= io_inputs_8;
    end else if (_T_14) begin
      _T_34 <= io_inputs_7;
    end else if (_T_12) begin
      _T_34 <= io_inputs_6;
    end else if (_T_10) begin
      _T_34 <= io_inputs_5;
    end else if (_T_8) begin
      _T_34 <= io_inputs_4;
    end else if (_T_6) begin
      _T_34 <= io_inputs_3;
    end else if (_T_4) begin
      _T_34 <= io_inputs_2;
    end else if (_T_2) begin
      _T_34 <= io_inputs_1;
    end else if (_T) begin
      _T_34 <= io_inputs_0;
    end else begin
      _T_34 <= 33'h0;
    end
  end
endmodule
module CfgMem_16(
  input          clock,
  input          reset,
  input          io_cfgEn,
  input  [3:0]   io_cfgAddr,
  input  [31:0]  io_cfgData,
  output [340:0] io_cfgOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  _T = io_cfgAddr == 4'h0; // @[CfgMem.scala 20:71]
  wire  _T_1 = io_cfgEn & _T; // @[CfgMem.scala 20:57]
  reg [31:0] outWire_0; // @[Reg.scala 27:20]
  wire  _T_3 = io_cfgAddr == 4'h1; // @[CfgMem.scala 20:71]
  wire  _T_4 = io_cfgEn & _T_3; // @[CfgMem.scala 20:57]
  reg [31:0] outWire_1; // @[Reg.scala 27:20]
  wire  _T_6 = io_cfgAddr == 4'h2; // @[CfgMem.scala 20:71]
  wire  _T_7 = io_cfgEn & _T_6; // @[CfgMem.scala 20:57]
  reg [31:0] outWire_2; // @[Reg.scala 27:20]
  wire  _T_9 = io_cfgAddr == 4'h3; // @[CfgMem.scala 20:71]
  wire  _T_10 = io_cfgEn & _T_9; // @[CfgMem.scala 20:57]
  reg [31:0] outWire_3; // @[Reg.scala 27:20]
  wire  _T_12 = io_cfgAddr == 4'h4; // @[CfgMem.scala 20:71]
  wire  _T_13 = io_cfgEn & _T_12; // @[CfgMem.scala 20:57]
  reg [31:0] outWire_4; // @[Reg.scala 27:20]
  wire  _T_15 = io_cfgAddr == 4'h5; // @[CfgMem.scala 20:71]
  wire  _T_16 = io_cfgEn & _T_15; // @[CfgMem.scala 20:57]
  reg [31:0] outWire_5; // @[Reg.scala 27:20]
  wire  _T_18 = io_cfgAddr == 4'h6; // @[CfgMem.scala 20:71]
  wire  _T_19 = io_cfgEn & _T_18; // @[CfgMem.scala 20:57]
  reg [31:0] outWire_6; // @[Reg.scala 27:20]
  wire  _T_21 = io_cfgAddr == 4'h7; // @[CfgMem.scala 20:71]
  wire  _T_22 = io_cfgEn & _T_21; // @[CfgMem.scala 20:57]
  reg [31:0] outWire_7; // @[Reg.scala 27:20]
  wire  _T_24 = io_cfgAddr == 4'h8; // @[CfgMem.scala 20:71]
  wire  _T_25 = io_cfgEn & _T_24; // @[CfgMem.scala 20:57]
  reg [31:0] outWire_8; // @[Reg.scala 27:20]
  wire  _T_27 = io_cfgAddr == 4'h9; // @[CfgMem.scala 20:71]
  wire  _T_28 = io_cfgEn & _T_27; // @[CfgMem.scala 20:57]
  reg [31:0] outWire_9; // @[Reg.scala 27:20]
  wire  _T_30 = io_cfgAddr == 4'ha; // @[CfgMem.scala 20:71]
  wire  _T_31 = io_cfgEn & _T_30; // @[CfgMem.scala 20:57]
  reg [31:0] outWire_10; // @[Reg.scala 27:20]
  wire [159:0] _T_36 = {outWire_4,outWire_3,outWire_2,outWire_1,outWire_0}; // @[Cat.scala 29:58]
  wire [351:0] _T_42 = {outWire_10,outWire_9,outWire_8,outWire_7,outWire_6,outWire_5,_T_36}; // @[Cat.scala 29:58]
  assign io_cfgOut = _T_42[340:0]; // @[CfgMem.scala 22:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  outWire_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  outWire_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  outWire_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  outWire_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  outWire_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  outWire_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  outWire_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  outWire_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  outWire_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  outWire_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  outWire_10 = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      outWire_0 <= 32'h0;
    end else if (_T_1) begin
      outWire_0 <= io_cfgData;
    end
    if (reset) begin
      outWire_1 <= 32'h0;
    end else if (_T_4) begin
      outWire_1 <= io_cfgData;
    end
    if (reset) begin
      outWire_2 <= 32'h0;
    end else if (_T_7) begin
      outWire_2 <= io_cfgData;
    end
    if (reset) begin
      outWire_3 <= 32'h0;
    end else if (_T_10) begin
      outWire_3 <= io_cfgData;
    end
    if (reset) begin
      outWire_4 <= 32'h0;
    end else if (_T_13) begin
      outWire_4 <= io_cfgData;
    end
    if (reset) begin
      outWire_5 <= 32'h0;
    end else if (_T_16) begin
      outWire_5 <= io_cfgData;
    end
    if (reset) begin
      outWire_6 <= 32'h0;
    end else if (_T_19) begin
      outWire_6 <= io_cfgData;
    end
    if (reset) begin
      outWire_7 <= 32'h0;
    end else if (_T_22) begin
      outWire_7 <= io_cfgData;
    end
    if (reset) begin
      outWire_8 <= 32'h0;
    end else if (_T_25) begin
      outWire_8 <= io_cfgData;
    end
    if (reset) begin
      outWire_9 <= 32'h0;
    end else if (_T_28) begin
      outWire_9 <= io_cfgData;
    end
    if (reset) begin
      outWire_10 <= 32'h0;
    end else if (_T_31) begin
      outWire_10 <= io_cfgData;
    end
  end
endmodule
module matrixFCdevice0(
  input         clock,
  input         reset,
  input         io_cfgEn,
  input  [3:0]  io_cfgAddr,
  input  [31:0] io_cfgData,
  input  [32:0] io_inputs_0,
  input  [32:0] io_inputs_1,
  input  [32:0] io_inputs_2,
  input  [32:0] io_inputs_3,
  input  [32:0] io_inputs_4,
  input  [32:0] io_inputs_5,
  input  [32:0] io_inputs_6,
  input  [32:0] io_inputs_7,
  input  [32:0] io_inputs_8,
  input  [32:0] io_inputs_9,
  input  [32:0] io_inputs_10,
  input  [32:0] io_inputs_11,
  input  [32:0] io_inputs_12,
  input  [32:0] io_inputs_13,
  input  [32:0] io_inputs_14,
  input  [32:0] io_inputs_15,
  input  [32:0] io_inputs_16,
  output [32:0] io_outputs_0,
  output [32:0] io_outputs_1,
  output [32:0] io_outputs_2,
  output [32:0] io_outputs_3,
  output [32:0] io_outputs_4,
  output [32:0] io_outputs_5,
  output [32:0] io_outputs_6,
  output [32:0] io_outputs_7,
  output [32:0] io_outputs_8,
  output [32:0] io_outputs_9,
  output [32:0] io_outputs_10,
  output [32:0] io_outputs_11,
  output [32:0] io_outputs_12,
  output [32:0] io_outputs_13,
  output [32:0] io_outputs_14,
  output [32:0] io_outputs_15,
  output [32:0] io_outputs_16
);
  wire [31:0] ConstUnit0_io_cfg; // @[TopModule.scala 192:48]
  wire [32:0] ConstUnit0_io_outputs_0; // @[TopModule.scala 192:48]
  wire [31:0] ConstUnit1_io_cfg; // @[TopModule.scala 192:48]
  wire [32:0] ConstUnit1_io_outputs_0; // @[TopModule.scala 192:48]
  wire [31:0] ConstUnit2_io_cfg; // @[TopModule.scala 192:48]
  wire [32:0] ConstUnit2_io_outputs_0; // @[TopModule.scala 192:48]
  wire [31:0] ConstUnit3_io_cfg; // @[TopModule.scala 192:48]
  wire [32:0] ConstUnit3_io_outputs_0; // @[TopModule.scala 192:48]
  wire [31:0] ConstUnit4_io_cfg; // @[TopModule.scala 192:48]
  wire [32:0] ConstUnit4_io_outputs_0; // @[TopModule.scala 192:48]
  wire [31:0] ConstUnit5_io_cfg; // @[TopModule.scala 192:48]
  wire [32:0] ConstUnit5_io_outputs_0; // @[TopModule.scala 192:48]
  wire [31:0] ConstUnit6_io_cfg; // @[TopModule.scala 192:48]
  wire [32:0] ConstUnit6_io_outputs_0; // @[TopModule.scala 192:48]
  wire [31:0] ConstUnit7_io_cfg; // @[TopModule.scala 192:48]
  wire [32:0] ConstUnit7_io_outputs_0; // @[TopModule.scala 192:48]
  wire [4:0] MUX0_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX1_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX2_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX3_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX4_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX5_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX6_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX7_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX8_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX9_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX10_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX11_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX12_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX13_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX14_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX15_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_outputs_0; // @[TopModule.scala 199:48]
  wire  MUXR0_clock; // @[TopModule.scala 205:48]
  wire  MUXR0_reset; // @[TopModule.scala 205:48]
  wire [4:0] MUXR0_io_cfg; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_0; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_1; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_2; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_3; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_4; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_5; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_6; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_7; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_8; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_9; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_10; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_11; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_12; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_13; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_14; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_15; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_16; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_outputs_0; // @[TopModule.scala 205:48]
  wire  CfgMem_clock; // @[TopModule.scala 232:29]
  wire  CfgMem_reset; // @[TopModule.scala 232:29]
  wire  CfgMem_io_cfgEn; // @[TopModule.scala 232:29]
  wire [3:0] CfgMem_io_cfgAddr; // @[TopModule.scala 232:29]
  wire [31:0] CfgMem_io_cfgData; // @[TopModule.scala 232:29]
  wire [340:0] CfgMem_io_cfgOut; // @[TopModule.scala 232:29]
  ConstUnit0 ConstUnit0 ( // @[TopModule.scala 192:48]
    .io_cfg(ConstUnit0_io_cfg),
    .io_outputs_0(ConstUnit0_io_outputs_0)
  );
  ConstUnit0 ConstUnit1 ( // @[TopModule.scala 192:48]
    .io_cfg(ConstUnit1_io_cfg),
    .io_outputs_0(ConstUnit1_io_outputs_0)
  );
  ConstUnit0 ConstUnit2 ( // @[TopModule.scala 192:48]
    .io_cfg(ConstUnit2_io_cfg),
    .io_outputs_0(ConstUnit2_io_outputs_0)
  );
  ConstUnit0 ConstUnit3 ( // @[TopModule.scala 192:48]
    .io_cfg(ConstUnit3_io_cfg),
    .io_outputs_0(ConstUnit3_io_outputs_0)
  );
  ConstUnit0 ConstUnit4 ( // @[TopModule.scala 192:48]
    .io_cfg(ConstUnit4_io_cfg),
    .io_outputs_0(ConstUnit4_io_outputs_0)
  );
  ConstUnit0 ConstUnit5 ( // @[TopModule.scala 192:48]
    .io_cfg(ConstUnit5_io_cfg),
    .io_outputs_0(ConstUnit5_io_outputs_0)
  );
  ConstUnit0 ConstUnit6 ( // @[TopModule.scala 192:48]
    .io_cfg(ConstUnit6_io_cfg),
    .io_outputs_0(ConstUnit6_io_outputs_0)
  );
  ConstUnit0 ConstUnit7 ( // @[TopModule.scala 192:48]
    .io_cfg(ConstUnit7_io_cfg),
    .io_outputs_0(ConstUnit7_io_outputs_0)
  );
  MUX0 MUX0 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX0_io_cfg),
    .io_inputs_0(MUX0_io_inputs_0),
    .io_inputs_1(MUX0_io_inputs_1),
    .io_inputs_2(MUX0_io_inputs_2),
    .io_inputs_3(MUX0_io_inputs_3),
    .io_inputs_4(MUX0_io_inputs_4),
    .io_inputs_5(MUX0_io_inputs_5),
    .io_inputs_6(MUX0_io_inputs_6),
    .io_inputs_7(MUX0_io_inputs_7),
    .io_inputs_8(MUX0_io_inputs_8),
    .io_inputs_9(MUX0_io_inputs_9),
    .io_inputs_10(MUX0_io_inputs_10),
    .io_inputs_11(MUX0_io_inputs_11),
    .io_inputs_12(MUX0_io_inputs_12),
    .io_inputs_13(MUX0_io_inputs_13),
    .io_inputs_14(MUX0_io_inputs_14),
    .io_inputs_15(MUX0_io_inputs_15),
    .io_inputs_16(MUX0_io_inputs_16),
    .io_outputs_0(MUX0_io_outputs_0)
  );
  MUX0 MUX1 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX1_io_cfg),
    .io_inputs_0(MUX1_io_inputs_0),
    .io_inputs_1(MUX1_io_inputs_1),
    .io_inputs_2(MUX1_io_inputs_2),
    .io_inputs_3(MUX1_io_inputs_3),
    .io_inputs_4(MUX1_io_inputs_4),
    .io_inputs_5(MUX1_io_inputs_5),
    .io_inputs_6(MUX1_io_inputs_6),
    .io_inputs_7(MUX1_io_inputs_7),
    .io_inputs_8(MUX1_io_inputs_8),
    .io_inputs_9(MUX1_io_inputs_9),
    .io_inputs_10(MUX1_io_inputs_10),
    .io_inputs_11(MUX1_io_inputs_11),
    .io_inputs_12(MUX1_io_inputs_12),
    .io_inputs_13(MUX1_io_inputs_13),
    .io_inputs_14(MUX1_io_inputs_14),
    .io_inputs_15(MUX1_io_inputs_15),
    .io_inputs_16(MUX1_io_inputs_16),
    .io_outputs_0(MUX1_io_outputs_0)
  );
  MUX0 MUX2 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX2_io_cfg),
    .io_inputs_0(MUX2_io_inputs_0),
    .io_inputs_1(MUX2_io_inputs_1),
    .io_inputs_2(MUX2_io_inputs_2),
    .io_inputs_3(MUX2_io_inputs_3),
    .io_inputs_4(MUX2_io_inputs_4),
    .io_inputs_5(MUX2_io_inputs_5),
    .io_inputs_6(MUX2_io_inputs_6),
    .io_inputs_7(MUX2_io_inputs_7),
    .io_inputs_8(MUX2_io_inputs_8),
    .io_inputs_9(MUX2_io_inputs_9),
    .io_inputs_10(MUX2_io_inputs_10),
    .io_inputs_11(MUX2_io_inputs_11),
    .io_inputs_12(MUX2_io_inputs_12),
    .io_inputs_13(MUX2_io_inputs_13),
    .io_inputs_14(MUX2_io_inputs_14),
    .io_inputs_15(MUX2_io_inputs_15),
    .io_inputs_16(MUX2_io_inputs_16),
    .io_outputs_0(MUX2_io_outputs_0)
  );
  MUX0 MUX3 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX3_io_cfg),
    .io_inputs_0(MUX3_io_inputs_0),
    .io_inputs_1(MUX3_io_inputs_1),
    .io_inputs_2(MUX3_io_inputs_2),
    .io_inputs_3(MUX3_io_inputs_3),
    .io_inputs_4(MUX3_io_inputs_4),
    .io_inputs_5(MUX3_io_inputs_5),
    .io_inputs_6(MUX3_io_inputs_6),
    .io_inputs_7(MUX3_io_inputs_7),
    .io_inputs_8(MUX3_io_inputs_8),
    .io_inputs_9(MUX3_io_inputs_9),
    .io_inputs_10(MUX3_io_inputs_10),
    .io_inputs_11(MUX3_io_inputs_11),
    .io_inputs_12(MUX3_io_inputs_12),
    .io_inputs_13(MUX3_io_inputs_13),
    .io_inputs_14(MUX3_io_inputs_14),
    .io_inputs_15(MUX3_io_inputs_15),
    .io_inputs_16(MUX3_io_inputs_16),
    .io_outputs_0(MUX3_io_outputs_0)
  );
  MUX0 MUX4 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX4_io_cfg),
    .io_inputs_0(MUX4_io_inputs_0),
    .io_inputs_1(MUX4_io_inputs_1),
    .io_inputs_2(MUX4_io_inputs_2),
    .io_inputs_3(MUX4_io_inputs_3),
    .io_inputs_4(MUX4_io_inputs_4),
    .io_inputs_5(MUX4_io_inputs_5),
    .io_inputs_6(MUX4_io_inputs_6),
    .io_inputs_7(MUX4_io_inputs_7),
    .io_inputs_8(MUX4_io_inputs_8),
    .io_inputs_9(MUX4_io_inputs_9),
    .io_inputs_10(MUX4_io_inputs_10),
    .io_inputs_11(MUX4_io_inputs_11),
    .io_inputs_12(MUX4_io_inputs_12),
    .io_inputs_13(MUX4_io_inputs_13),
    .io_inputs_14(MUX4_io_inputs_14),
    .io_inputs_15(MUX4_io_inputs_15),
    .io_inputs_16(MUX4_io_inputs_16),
    .io_outputs_0(MUX4_io_outputs_0)
  );
  MUX0 MUX5 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX5_io_cfg),
    .io_inputs_0(MUX5_io_inputs_0),
    .io_inputs_1(MUX5_io_inputs_1),
    .io_inputs_2(MUX5_io_inputs_2),
    .io_inputs_3(MUX5_io_inputs_3),
    .io_inputs_4(MUX5_io_inputs_4),
    .io_inputs_5(MUX5_io_inputs_5),
    .io_inputs_6(MUX5_io_inputs_6),
    .io_inputs_7(MUX5_io_inputs_7),
    .io_inputs_8(MUX5_io_inputs_8),
    .io_inputs_9(MUX5_io_inputs_9),
    .io_inputs_10(MUX5_io_inputs_10),
    .io_inputs_11(MUX5_io_inputs_11),
    .io_inputs_12(MUX5_io_inputs_12),
    .io_inputs_13(MUX5_io_inputs_13),
    .io_inputs_14(MUX5_io_inputs_14),
    .io_inputs_15(MUX5_io_inputs_15),
    .io_inputs_16(MUX5_io_inputs_16),
    .io_outputs_0(MUX5_io_outputs_0)
  );
  MUX0 MUX6 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX6_io_cfg),
    .io_inputs_0(MUX6_io_inputs_0),
    .io_inputs_1(MUX6_io_inputs_1),
    .io_inputs_2(MUX6_io_inputs_2),
    .io_inputs_3(MUX6_io_inputs_3),
    .io_inputs_4(MUX6_io_inputs_4),
    .io_inputs_5(MUX6_io_inputs_5),
    .io_inputs_6(MUX6_io_inputs_6),
    .io_inputs_7(MUX6_io_inputs_7),
    .io_inputs_8(MUX6_io_inputs_8),
    .io_inputs_9(MUX6_io_inputs_9),
    .io_inputs_10(MUX6_io_inputs_10),
    .io_inputs_11(MUX6_io_inputs_11),
    .io_inputs_12(MUX6_io_inputs_12),
    .io_inputs_13(MUX6_io_inputs_13),
    .io_inputs_14(MUX6_io_inputs_14),
    .io_inputs_15(MUX6_io_inputs_15),
    .io_inputs_16(MUX6_io_inputs_16),
    .io_outputs_0(MUX6_io_outputs_0)
  );
  MUX0 MUX7 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX7_io_cfg),
    .io_inputs_0(MUX7_io_inputs_0),
    .io_inputs_1(MUX7_io_inputs_1),
    .io_inputs_2(MUX7_io_inputs_2),
    .io_inputs_3(MUX7_io_inputs_3),
    .io_inputs_4(MUX7_io_inputs_4),
    .io_inputs_5(MUX7_io_inputs_5),
    .io_inputs_6(MUX7_io_inputs_6),
    .io_inputs_7(MUX7_io_inputs_7),
    .io_inputs_8(MUX7_io_inputs_8),
    .io_inputs_9(MUX7_io_inputs_9),
    .io_inputs_10(MUX7_io_inputs_10),
    .io_inputs_11(MUX7_io_inputs_11),
    .io_inputs_12(MUX7_io_inputs_12),
    .io_inputs_13(MUX7_io_inputs_13),
    .io_inputs_14(MUX7_io_inputs_14),
    .io_inputs_15(MUX7_io_inputs_15),
    .io_inputs_16(MUX7_io_inputs_16),
    .io_outputs_0(MUX7_io_outputs_0)
  );
  MUX8 MUX8 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX8_io_cfg),
    .io_inputs_0(MUX8_io_inputs_0),
    .io_inputs_1(MUX8_io_inputs_1),
    .io_inputs_2(MUX8_io_inputs_2),
    .io_inputs_3(MUX8_io_inputs_3),
    .io_inputs_4(MUX8_io_inputs_4),
    .io_inputs_5(MUX8_io_inputs_5),
    .io_inputs_6(MUX8_io_inputs_6),
    .io_inputs_7(MUX8_io_inputs_7),
    .io_inputs_8(MUX8_io_inputs_8),
    .io_inputs_9(MUX8_io_inputs_9),
    .io_inputs_10(MUX8_io_inputs_10),
    .io_inputs_11(MUX8_io_inputs_11),
    .io_inputs_12(MUX8_io_inputs_12),
    .io_inputs_13(MUX8_io_inputs_13),
    .io_inputs_14(MUX8_io_inputs_14),
    .io_inputs_15(MUX8_io_inputs_15),
    .io_inputs_16(MUX8_io_inputs_16),
    .io_inputs_17(MUX8_io_inputs_17),
    .io_outputs_0(MUX8_io_outputs_0)
  );
  MUX8 MUX9 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX9_io_cfg),
    .io_inputs_0(MUX9_io_inputs_0),
    .io_inputs_1(MUX9_io_inputs_1),
    .io_inputs_2(MUX9_io_inputs_2),
    .io_inputs_3(MUX9_io_inputs_3),
    .io_inputs_4(MUX9_io_inputs_4),
    .io_inputs_5(MUX9_io_inputs_5),
    .io_inputs_6(MUX9_io_inputs_6),
    .io_inputs_7(MUX9_io_inputs_7),
    .io_inputs_8(MUX9_io_inputs_8),
    .io_inputs_9(MUX9_io_inputs_9),
    .io_inputs_10(MUX9_io_inputs_10),
    .io_inputs_11(MUX9_io_inputs_11),
    .io_inputs_12(MUX9_io_inputs_12),
    .io_inputs_13(MUX9_io_inputs_13),
    .io_inputs_14(MUX9_io_inputs_14),
    .io_inputs_15(MUX9_io_inputs_15),
    .io_inputs_16(MUX9_io_inputs_16),
    .io_inputs_17(MUX9_io_inputs_17),
    .io_outputs_0(MUX9_io_outputs_0)
  );
  MUX8 MUX10 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX10_io_cfg),
    .io_inputs_0(MUX10_io_inputs_0),
    .io_inputs_1(MUX10_io_inputs_1),
    .io_inputs_2(MUX10_io_inputs_2),
    .io_inputs_3(MUX10_io_inputs_3),
    .io_inputs_4(MUX10_io_inputs_4),
    .io_inputs_5(MUX10_io_inputs_5),
    .io_inputs_6(MUX10_io_inputs_6),
    .io_inputs_7(MUX10_io_inputs_7),
    .io_inputs_8(MUX10_io_inputs_8),
    .io_inputs_9(MUX10_io_inputs_9),
    .io_inputs_10(MUX10_io_inputs_10),
    .io_inputs_11(MUX10_io_inputs_11),
    .io_inputs_12(MUX10_io_inputs_12),
    .io_inputs_13(MUX10_io_inputs_13),
    .io_inputs_14(MUX10_io_inputs_14),
    .io_inputs_15(MUX10_io_inputs_15),
    .io_inputs_16(MUX10_io_inputs_16),
    .io_inputs_17(MUX10_io_inputs_17),
    .io_outputs_0(MUX10_io_outputs_0)
  );
  MUX8 MUX11 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX11_io_cfg),
    .io_inputs_0(MUX11_io_inputs_0),
    .io_inputs_1(MUX11_io_inputs_1),
    .io_inputs_2(MUX11_io_inputs_2),
    .io_inputs_3(MUX11_io_inputs_3),
    .io_inputs_4(MUX11_io_inputs_4),
    .io_inputs_5(MUX11_io_inputs_5),
    .io_inputs_6(MUX11_io_inputs_6),
    .io_inputs_7(MUX11_io_inputs_7),
    .io_inputs_8(MUX11_io_inputs_8),
    .io_inputs_9(MUX11_io_inputs_9),
    .io_inputs_10(MUX11_io_inputs_10),
    .io_inputs_11(MUX11_io_inputs_11),
    .io_inputs_12(MUX11_io_inputs_12),
    .io_inputs_13(MUX11_io_inputs_13),
    .io_inputs_14(MUX11_io_inputs_14),
    .io_inputs_15(MUX11_io_inputs_15),
    .io_inputs_16(MUX11_io_inputs_16),
    .io_inputs_17(MUX11_io_inputs_17),
    .io_outputs_0(MUX11_io_outputs_0)
  );
  MUX8 MUX12 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX12_io_cfg),
    .io_inputs_0(MUX12_io_inputs_0),
    .io_inputs_1(MUX12_io_inputs_1),
    .io_inputs_2(MUX12_io_inputs_2),
    .io_inputs_3(MUX12_io_inputs_3),
    .io_inputs_4(MUX12_io_inputs_4),
    .io_inputs_5(MUX12_io_inputs_5),
    .io_inputs_6(MUX12_io_inputs_6),
    .io_inputs_7(MUX12_io_inputs_7),
    .io_inputs_8(MUX12_io_inputs_8),
    .io_inputs_9(MUX12_io_inputs_9),
    .io_inputs_10(MUX12_io_inputs_10),
    .io_inputs_11(MUX12_io_inputs_11),
    .io_inputs_12(MUX12_io_inputs_12),
    .io_inputs_13(MUX12_io_inputs_13),
    .io_inputs_14(MUX12_io_inputs_14),
    .io_inputs_15(MUX12_io_inputs_15),
    .io_inputs_16(MUX12_io_inputs_16),
    .io_inputs_17(MUX12_io_inputs_17),
    .io_outputs_0(MUX12_io_outputs_0)
  );
  MUX8 MUX13 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX13_io_cfg),
    .io_inputs_0(MUX13_io_inputs_0),
    .io_inputs_1(MUX13_io_inputs_1),
    .io_inputs_2(MUX13_io_inputs_2),
    .io_inputs_3(MUX13_io_inputs_3),
    .io_inputs_4(MUX13_io_inputs_4),
    .io_inputs_5(MUX13_io_inputs_5),
    .io_inputs_6(MUX13_io_inputs_6),
    .io_inputs_7(MUX13_io_inputs_7),
    .io_inputs_8(MUX13_io_inputs_8),
    .io_inputs_9(MUX13_io_inputs_9),
    .io_inputs_10(MUX13_io_inputs_10),
    .io_inputs_11(MUX13_io_inputs_11),
    .io_inputs_12(MUX13_io_inputs_12),
    .io_inputs_13(MUX13_io_inputs_13),
    .io_inputs_14(MUX13_io_inputs_14),
    .io_inputs_15(MUX13_io_inputs_15),
    .io_inputs_16(MUX13_io_inputs_16),
    .io_inputs_17(MUX13_io_inputs_17),
    .io_outputs_0(MUX13_io_outputs_0)
  );
  MUX8 MUX14 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX14_io_cfg),
    .io_inputs_0(MUX14_io_inputs_0),
    .io_inputs_1(MUX14_io_inputs_1),
    .io_inputs_2(MUX14_io_inputs_2),
    .io_inputs_3(MUX14_io_inputs_3),
    .io_inputs_4(MUX14_io_inputs_4),
    .io_inputs_5(MUX14_io_inputs_5),
    .io_inputs_6(MUX14_io_inputs_6),
    .io_inputs_7(MUX14_io_inputs_7),
    .io_inputs_8(MUX14_io_inputs_8),
    .io_inputs_9(MUX14_io_inputs_9),
    .io_inputs_10(MUX14_io_inputs_10),
    .io_inputs_11(MUX14_io_inputs_11),
    .io_inputs_12(MUX14_io_inputs_12),
    .io_inputs_13(MUX14_io_inputs_13),
    .io_inputs_14(MUX14_io_inputs_14),
    .io_inputs_15(MUX14_io_inputs_15),
    .io_inputs_16(MUX14_io_inputs_16),
    .io_inputs_17(MUX14_io_inputs_17),
    .io_outputs_0(MUX14_io_outputs_0)
  );
  MUX8 MUX15 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX15_io_cfg),
    .io_inputs_0(MUX15_io_inputs_0),
    .io_inputs_1(MUX15_io_inputs_1),
    .io_inputs_2(MUX15_io_inputs_2),
    .io_inputs_3(MUX15_io_inputs_3),
    .io_inputs_4(MUX15_io_inputs_4),
    .io_inputs_5(MUX15_io_inputs_5),
    .io_inputs_6(MUX15_io_inputs_6),
    .io_inputs_7(MUX15_io_inputs_7),
    .io_inputs_8(MUX15_io_inputs_8),
    .io_inputs_9(MUX15_io_inputs_9),
    .io_inputs_10(MUX15_io_inputs_10),
    .io_inputs_11(MUX15_io_inputs_11),
    .io_inputs_12(MUX15_io_inputs_12),
    .io_inputs_13(MUX15_io_inputs_13),
    .io_inputs_14(MUX15_io_inputs_14),
    .io_inputs_15(MUX15_io_inputs_15),
    .io_inputs_16(MUX15_io_inputs_16),
    .io_inputs_17(MUX15_io_inputs_17),
    .io_outputs_0(MUX15_io_outputs_0)
  );
  MUXR0 MUXR0 ( // @[TopModule.scala 205:48]
    .clock(MUXR0_clock),
    .reset(MUXR0_reset),
    .io_cfg(MUXR0_io_cfg),
    .io_inputs_0(MUXR0_io_inputs_0),
    .io_inputs_1(MUXR0_io_inputs_1),
    .io_inputs_2(MUXR0_io_inputs_2),
    .io_inputs_3(MUXR0_io_inputs_3),
    .io_inputs_4(MUXR0_io_inputs_4),
    .io_inputs_5(MUXR0_io_inputs_5),
    .io_inputs_6(MUXR0_io_inputs_6),
    .io_inputs_7(MUXR0_io_inputs_7),
    .io_inputs_8(MUXR0_io_inputs_8),
    .io_inputs_9(MUXR0_io_inputs_9),
    .io_inputs_10(MUXR0_io_inputs_10),
    .io_inputs_11(MUXR0_io_inputs_11),
    .io_inputs_12(MUXR0_io_inputs_12),
    .io_inputs_13(MUXR0_io_inputs_13),
    .io_inputs_14(MUXR0_io_inputs_14),
    .io_inputs_15(MUXR0_io_inputs_15),
    .io_inputs_16(MUXR0_io_inputs_16),
    .io_outputs_0(MUXR0_io_outputs_0)
  );
  CfgMem_16 CfgMem ( // @[TopModule.scala 232:29]
    .clock(CfgMem_clock),
    .reset(CfgMem_reset),
    .io_cfgEn(CfgMem_io_cfgEn),
    .io_cfgAddr(CfgMem_io_cfgAddr),
    .io_cfgData(CfgMem_io_cfgData),
    .io_cfgOut(CfgMem_io_cfgOut)
  );
  assign io_outputs_0 = MUXR0_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_1 = MUX0_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_2 = MUX1_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_3 = MUX2_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_4 = MUX3_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_5 = MUX4_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_6 = MUX5_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_7 = MUX6_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_8 = MUX7_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_9 = MUX8_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_10 = MUX9_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_11 = MUX10_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_12 = MUX11_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_13 = MUX12_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_14 = MUX13_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_15 = MUX14_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_16 = MUX15_io_outputs_0; // @[TopModule.scala 392:22]
  assign ConstUnit0_io_cfg = CfgMem_io_cfgOut[31:0]; // @[TopModule.scala 259:94]
  assign ConstUnit1_io_cfg = CfgMem_io_cfgOut[63:32]; // @[TopModule.scala 259:94]
  assign ConstUnit2_io_cfg = CfgMem_io_cfgOut[95:64]; // @[TopModule.scala 259:94]
  assign ConstUnit3_io_cfg = CfgMem_io_cfgOut[127:96]; // @[TopModule.scala 259:94]
  assign ConstUnit4_io_cfg = CfgMem_io_cfgOut[159:128]; // @[TopModule.scala 259:94]
  assign ConstUnit5_io_cfg = CfgMem_io_cfgOut[191:160]; // @[TopModule.scala 259:94]
  assign ConstUnit6_io_cfg = CfgMem_io_cfgOut[223:192]; // @[TopModule.scala 259:94]
  assign ConstUnit7_io_cfg = CfgMem_io_cfgOut[255:224]; // @[TopModule.scala 259:94]
  assign MUX0_io_cfg = CfgMem_io_cfgOut[260:256]; // @[TopModule.scala 261:98]
  assign MUX0_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX1_io_cfg = CfgMem_io_cfgOut[265:261]; // @[TopModule.scala 261:98]
  assign MUX1_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX2_io_cfg = CfgMem_io_cfgOut[270:266]; // @[TopModule.scala 261:98]
  assign MUX2_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX3_io_cfg = CfgMem_io_cfgOut[275:271]; // @[TopModule.scala 261:98]
  assign MUX3_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX4_io_cfg = CfgMem_io_cfgOut[280:276]; // @[TopModule.scala 261:98]
  assign MUX4_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX5_io_cfg = CfgMem_io_cfgOut[285:281]; // @[TopModule.scala 261:98]
  assign MUX5_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX6_io_cfg = CfgMem_io_cfgOut[290:286]; // @[TopModule.scala 261:98]
  assign MUX6_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX7_io_cfg = CfgMem_io_cfgOut[295:291]; // @[TopModule.scala 261:98]
  assign MUX7_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX8_io_cfg = CfgMem_io_cfgOut[300:296]; // @[TopModule.scala 261:98]
  assign MUX8_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_17 = ConstUnit0_io_outputs_0; // @[TopModule.scala 392:22]
  assign MUX9_io_cfg = CfgMem_io_cfgOut[305:301]; // @[TopModule.scala 261:98]
  assign MUX9_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_17 = ConstUnit1_io_outputs_0; // @[TopModule.scala 392:22]
  assign MUX10_io_cfg = CfgMem_io_cfgOut[310:306]; // @[TopModule.scala 261:98]
  assign MUX10_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_17 = ConstUnit2_io_outputs_0; // @[TopModule.scala 392:22]
  assign MUX11_io_cfg = CfgMem_io_cfgOut[315:311]; // @[TopModule.scala 261:98]
  assign MUX11_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_17 = ConstUnit3_io_outputs_0; // @[TopModule.scala 392:22]
  assign MUX12_io_cfg = CfgMem_io_cfgOut[320:316]; // @[TopModule.scala 261:98]
  assign MUX12_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_17 = ConstUnit4_io_outputs_0; // @[TopModule.scala 392:22]
  assign MUX13_io_cfg = CfgMem_io_cfgOut[325:321]; // @[TopModule.scala 261:98]
  assign MUX13_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_17 = ConstUnit5_io_outputs_0; // @[TopModule.scala 392:22]
  assign MUX14_io_cfg = CfgMem_io_cfgOut[330:326]; // @[TopModule.scala 261:98]
  assign MUX14_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_17 = ConstUnit6_io_outputs_0; // @[TopModule.scala 392:22]
  assign MUX15_io_cfg = CfgMem_io_cfgOut[335:331]; // @[TopModule.scala 261:98]
  assign MUX15_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_17 = ConstUnit7_io_outputs_0; // @[TopModule.scala 392:22]
  assign MUXR0_clock = clock;
  assign MUXR0_reset = reset;
  assign MUXR0_io_cfg = CfgMem_io_cfgOut[340:336]; // @[TopModule.scala 262:100]
  assign MUXR0_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign CfgMem_clock = clock;
  assign CfgMem_reset = reset;
  assign CfgMem_io_cfgEn = io_cfgEn; // @[TopModule.scala 239:34]
  assign CfgMem_io_cfgAddr = io_cfgAddr; // @[TopModule.scala 244:30]
  assign CfgMem_io_cfgData = io_cfgData; // @[TopModule.scala 248:28]
endmodule
module MUX0_1(
  input  [4:0]  io_cfg,
  input  [32:0] io_inputs_0,
  input  [32:0] io_inputs_1,
  input  [32:0] io_inputs_2,
  input  [32:0] io_inputs_3,
  input  [32:0] io_inputs_4,
  input  [32:0] io_inputs_5,
  input  [32:0] io_inputs_6,
  input  [32:0] io_inputs_7,
  input  [32:0] io_inputs_8,
  input  [32:0] io_inputs_9,
  input  [32:0] io_inputs_10,
  input  [32:0] io_inputs_11,
  input  [32:0] io_inputs_12,
  input  [32:0] io_inputs_13,
  input  [32:0] io_inputs_14,
  input  [32:0] io_inputs_15,
  input  [32:0] io_inputs_16,
  input  [32:0] io_inputs_17,
  input  [32:0] io_inputs_18,
  input  [32:0] io_inputs_19,
  input  [32:0] io_inputs_20,
  input  [32:0] io_inputs_21,
  input  [32:0] io_inputs_22,
  input  [32:0] io_inputs_23,
  output [32:0] io_outputs_0
);
  wire  _T = 5'h0 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_1 = _T ? io_inputs_0 : 33'h0; // @[Mux.scala 80:57]
  wire  _T_2 = 5'h1 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_3 = _T_2 ? io_inputs_1 : _T_1; // @[Mux.scala 80:57]
  wire  _T_4 = 5'h2 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_5 = _T_4 ? io_inputs_2 : _T_3; // @[Mux.scala 80:57]
  wire  _T_6 = 5'h3 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_7 = _T_6 ? io_inputs_3 : _T_5; // @[Mux.scala 80:57]
  wire  _T_8 = 5'h4 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_9 = _T_8 ? io_inputs_4 : _T_7; // @[Mux.scala 80:57]
  wire  _T_10 = 5'h5 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_11 = _T_10 ? io_inputs_5 : _T_9; // @[Mux.scala 80:57]
  wire  _T_12 = 5'h6 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_13 = _T_12 ? io_inputs_6 : _T_11; // @[Mux.scala 80:57]
  wire  _T_14 = 5'h7 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_15 = _T_14 ? io_inputs_7 : _T_13; // @[Mux.scala 80:57]
  wire  _T_16 = 5'h8 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_17 = _T_16 ? io_inputs_8 : _T_15; // @[Mux.scala 80:57]
  wire  _T_18 = 5'h9 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_19 = _T_18 ? io_inputs_9 : _T_17; // @[Mux.scala 80:57]
  wire  _T_20 = 5'ha == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_21 = _T_20 ? io_inputs_10 : _T_19; // @[Mux.scala 80:57]
  wire  _T_22 = 5'hb == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_23 = _T_22 ? io_inputs_11 : _T_21; // @[Mux.scala 80:57]
  wire  _T_24 = 5'hc == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_25 = _T_24 ? io_inputs_12 : _T_23; // @[Mux.scala 80:57]
  wire  _T_26 = 5'hd == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_27 = _T_26 ? io_inputs_13 : _T_25; // @[Mux.scala 80:57]
  wire  _T_28 = 5'he == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_29 = _T_28 ? io_inputs_14 : _T_27; // @[Mux.scala 80:57]
  wire  _T_30 = 5'hf == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_31 = _T_30 ? io_inputs_15 : _T_29; // @[Mux.scala 80:57]
  wire  _T_32 = 5'h10 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_33 = _T_32 ? io_inputs_16 : _T_31; // @[Mux.scala 80:57]
  wire  _T_34 = 5'h11 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_35 = _T_34 ? io_inputs_17 : _T_33; // @[Mux.scala 80:57]
  wire  _T_36 = 5'h12 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_37 = _T_36 ? io_inputs_18 : _T_35; // @[Mux.scala 80:57]
  wire  _T_38 = 5'h13 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_39 = _T_38 ? io_inputs_19 : _T_37; // @[Mux.scala 80:57]
  wire  _T_40 = 5'h14 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_41 = _T_40 ? io_inputs_20 : _T_39; // @[Mux.scala 80:57]
  wire  _T_42 = 5'h15 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_43 = _T_42 ? io_inputs_21 : _T_41; // @[Mux.scala 80:57]
  wire  _T_44 = 5'h16 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_45 = _T_44 ? io_inputs_22 : _T_43; // @[Mux.scala 80:57]
  wire  _T_46 = 5'h17 == io_cfg; // @[Mux.scala 80:60]
  assign io_outputs_0 = _T_46 ? io_inputs_23 : _T_45; // @[Multiplexer.scala 16:17]
endmodule
module MUX8_1(
  input  [4:0]  io_cfg,
  input  [32:0] io_inputs_0,
  input  [32:0] io_inputs_1,
  input  [32:0] io_inputs_2,
  input  [32:0] io_inputs_3,
  input  [32:0] io_inputs_4,
  input  [32:0] io_inputs_5,
  input  [32:0] io_inputs_6,
  input  [32:0] io_inputs_7,
  input  [32:0] io_inputs_8,
  input  [32:0] io_inputs_9,
  input  [32:0] io_inputs_10,
  input  [32:0] io_inputs_11,
  input  [32:0] io_inputs_12,
  input  [32:0] io_inputs_13,
  input  [32:0] io_inputs_14,
  input  [32:0] io_inputs_15,
  input  [32:0] io_inputs_16,
  input  [32:0] io_inputs_17,
  input  [32:0] io_inputs_18,
  input  [32:0] io_inputs_19,
  input  [32:0] io_inputs_20,
  input  [32:0] io_inputs_21,
  input  [32:0] io_inputs_22,
  input  [32:0] io_inputs_23,
  input  [32:0] io_inputs_24,
  output [32:0] io_outputs_0
);
  wire  _T = 5'h0 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_1 = _T ? io_inputs_0 : 33'h0; // @[Mux.scala 80:57]
  wire  _T_2 = 5'h1 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_3 = _T_2 ? io_inputs_1 : _T_1; // @[Mux.scala 80:57]
  wire  _T_4 = 5'h2 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_5 = _T_4 ? io_inputs_2 : _T_3; // @[Mux.scala 80:57]
  wire  _T_6 = 5'h3 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_7 = _T_6 ? io_inputs_3 : _T_5; // @[Mux.scala 80:57]
  wire  _T_8 = 5'h4 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_9 = _T_8 ? io_inputs_4 : _T_7; // @[Mux.scala 80:57]
  wire  _T_10 = 5'h5 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_11 = _T_10 ? io_inputs_5 : _T_9; // @[Mux.scala 80:57]
  wire  _T_12 = 5'h6 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_13 = _T_12 ? io_inputs_6 : _T_11; // @[Mux.scala 80:57]
  wire  _T_14 = 5'h7 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_15 = _T_14 ? io_inputs_7 : _T_13; // @[Mux.scala 80:57]
  wire  _T_16 = 5'h8 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_17 = _T_16 ? io_inputs_8 : _T_15; // @[Mux.scala 80:57]
  wire  _T_18 = 5'h9 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_19 = _T_18 ? io_inputs_9 : _T_17; // @[Mux.scala 80:57]
  wire  _T_20 = 5'ha == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_21 = _T_20 ? io_inputs_10 : _T_19; // @[Mux.scala 80:57]
  wire  _T_22 = 5'hb == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_23 = _T_22 ? io_inputs_11 : _T_21; // @[Mux.scala 80:57]
  wire  _T_24 = 5'hc == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_25 = _T_24 ? io_inputs_12 : _T_23; // @[Mux.scala 80:57]
  wire  _T_26 = 5'hd == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_27 = _T_26 ? io_inputs_13 : _T_25; // @[Mux.scala 80:57]
  wire  _T_28 = 5'he == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_29 = _T_28 ? io_inputs_14 : _T_27; // @[Mux.scala 80:57]
  wire  _T_30 = 5'hf == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_31 = _T_30 ? io_inputs_15 : _T_29; // @[Mux.scala 80:57]
  wire  _T_32 = 5'h10 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_33 = _T_32 ? io_inputs_16 : _T_31; // @[Mux.scala 80:57]
  wire  _T_34 = 5'h11 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_35 = _T_34 ? io_inputs_17 : _T_33; // @[Mux.scala 80:57]
  wire  _T_36 = 5'h12 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_37 = _T_36 ? io_inputs_18 : _T_35; // @[Mux.scala 80:57]
  wire  _T_38 = 5'h13 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_39 = _T_38 ? io_inputs_19 : _T_37; // @[Mux.scala 80:57]
  wire  _T_40 = 5'h14 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_41 = _T_40 ? io_inputs_20 : _T_39; // @[Mux.scala 80:57]
  wire  _T_42 = 5'h15 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_43 = _T_42 ? io_inputs_21 : _T_41; // @[Mux.scala 80:57]
  wire  _T_44 = 5'h16 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_45 = _T_44 ? io_inputs_22 : _T_43; // @[Mux.scala 80:57]
  wire  _T_46 = 5'h17 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_47 = _T_46 ? io_inputs_23 : _T_45; // @[Mux.scala 80:57]
  wire  _T_48 = 5'h18 == io_cfg; // @[Mux.scala 80:60]
  assign io_outputs_0 = _T_48 ? io_inputs_24 : _T_47; // @[Multiplexer.scala 16:17]
endmodule
module MUXR0_1(
  input         clock,
  input         reset,
  input  [4:0]  io_cfg,
  input  [32:0] io_inputs_0,
  input  [32:0] io_inputs_1,
  input  [32:0] io_inputs_2,
  input  [32:0] io_inputs_3,
  input  [32:0] io_inputs_4,
  input  [32:0] io_inputs_5,
  input  [32:0] io_inputs_6,
  input  [32:0] io_inputs_7,
  input  [32:0] io_inputs_8,
  input  [32:0] io_inputs_9,
  input  [32:0] io_inputs_10,
  input  [32:0] io_inputs_11,
  input  [32:0] io_inputs_12,
  input  [32:0] io_inputs_13,
  input  [32:0] io_inputs_14,
  input  [32:0] io_inputs_15,
  input  [32:0] io_inputs_16,
  input  [32:0] io_inputs_17,
  input  [32:0] io_inputs_18,
  input  [32:0] io_inputs_19,
  input  [32:0] io_inputs_20,
  input  [32:0] io_inputs_21,
  input  [32:0] io_inputs_22,
  input  [32:0] io_inputs_23,
  output [32:0] io_outputs_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _T = 5'h0 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_2 = 5'h1 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_4 = 5'h2 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_6 = 5'h3 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_8 = 5'h4 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_10 = 5'h5 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_12 = 5'h6 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_14 = 5'h7 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_16 = 5'h8 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_18 = 5'h9 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_20 = 5'ha == io_cfg; // @[Mux.scala 80:60]
  wire  _T_22 = 5'hb == io_cfg; // @[Mux.scala 80:60]
  wire  _T_24 = 5'hc == io_cfg; // @[Mux.scala 80:60]
  wire  _T_26 = 5'hd == io_cfg; // @[Mux.scala 80:60]
  wire  _T_28 = 5'he == io_cfg; // @[Mux.scala 80:60]
  wire  _T_30 = 5'hf == io_cfg; // @[Mux.scala 80:60]
  wire  _T_32 = 5'h10 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_34 = 5'h11 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_36 = 5'h12 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_38 = 5'h13 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_40 = 5'h14 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_42 = 5'h15 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_44 = 5'h16 == io_cfg; // @[Mux.scala 80:60]
  wire  _T_46 = 5'h17 == io_cfg; // @[Mux.scala 80:60]
  reg [32:0] _T_48; // @[MultiplexerR.scala 16:27]
  assign io_outputs_0 = _T_48; // @[MultiplexerR.scala 16:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_48 = _RAND_0[32:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_48 <= 33'h0;
    end else if (_T_46) begin
      _T_48 <= io_inputs_23;
    end else if (_T_44) begin
      _T_48 <= io_inputs_22;
    end else if (_T_42) begin
      _T_48 <= io_inputs_21;
    end else if (_T_40) begin
      _T_48 <= io_inputs_20;
    end else if (_T_38) begin
      _T_48 <= io_inputs_19;
    end else if (_T_36) begin
      _T_48 <= io_inputs_18;
    end else if (_T_34) begin
      _T_48 <= io_inputs_17;
    end else if (_T_32) begin
      _T_48 <= io_inputs_16;
    end else if (_T_30) begin
      _T_48 <= io_inputs_15;
    end else if (_T_28) begin
      _T_48 <= io_inputs_14;
    end else if (_T_26) begin
      _T_48 <= io_inputs_13;
    end else if (_T_24) begin
      _T_48 <= io_inputs_12;
    end else if (_T_22) begin
      _T_48 <= io_inputs_11;
    end else if (_T_20) begin
      _T_48 <= io_inputs_10;
    end else if (_T_18) begin
      _T_48 <= io_inputs_9;
    end else if (_T_16) begin
      _T_48 <= io_inputs_8;
    end else if (_T_14) begin
      _T_48 <= io_inputs_7;
    end else if (_T_12) begin
      _T_48 <= io_inputs_6;
    end else if (_T_10) begin
      _T_48 <= io_inputs_5;
    end else if (_T_8) begin
      _T_48 <= io_inputs_4;
    end else if (_T_6) begin
      _T_48 <= io_inputs_3;
    end else if (_T_4) begin
      _T_48 <= io_inputs_2;
    end else if (_T_2) begin
      _T_48 <= io_inputs_1;
    end else if (_T) begin
      _T_48 <= io_inputs_0;
    end else begin
      _T_48 <= 33'h0;
    end
  end
endmodule
module matrixFCdevice1(
  input         clock,
  input         reset,
  input         io_cfgEn,
  input  [3:0]  io_cfgAddr,
  input  [31:0] io_cfgData,
  input  [32:0] io_inputs_0,
  input  [32:0] io_inputs_1,
  input  [32:0] io_inputs_2,
  input  [32:0] io_inputs_3,
  input  [32:0] io_inputs_4,
  input  [32:0] io_inputs_5,
  input  [32:0] io_inputs_6,
  input  [32:0] io_inputs_7,
  input  [32:0] io_inputs_8,
  input  [32:0] io_inputs_9,
  input  [32:0] io_inputs_10,
  input  [32:0] io_inputs_11,
  input  [32:0] io_inputs_12,
  input  [32:0] io_inputs_13,
  input  [32:0] io_inputs_14,
  input  [32:0] io_inputs_15,
  input  [32:0] io_inputs_16,
  input  [32:0] io_inputs_17,
  input  [32:0] io_inputs_18,
  input  [32:0] io_inputs_19,
  input  [32:0] io_inputs_20,
  input  [32:0] io_inputs_21,
  input  [32:0] io_inputs_22,
  input  [32:0] io_inputs_23,
  output [32:0] io_outputs_0,
  output [32:0] io_outputs_1,
  output [32:0] io_outputs_2,
  output [32:0] io_outputs_3,
  output [32:0] io_outputs_4,
  output [32:0] io_outputs_5,
  output [32:0] io_outputs_6,
  output [32:0] io_outputs_7,
  output [32:0] io_outputs_8,
  output [32:0] io_outputs_9,
  output [32:0] io_outputs_10,
  output [32:0] io_outputs_11,
  output [32:0] io_outputs_12,
  output [32:0] io_outputs_13,
  output [32:0] io_outputs_14,
  output [32:0] io_outputs_15,
  output [32:0] io_outputs_16
);
  wire [31:0] ConstUnit0_io_cfg; // @[TopModule.scala 192:48]
  wire [32:0] ConstUnit0_io_outputs_0; // @[TopModule.scala 192:48]
  wire [31:0] ConstUnit1_io_cfg; // @[TopModule.scala 192:48]
  wire [32:0] ConstUnit1_io_outputs_0; // @[TopModule.scala 192:48]
  wire [31:0] ConstUnit2_io_cfg; // @[TopModule.scala 192:48]
  wire [32:0] ConstUnit2_io_outputs_0; // @[TopModule.scala 192:48]
  wire [31:0] ConstUnit3_io_cfg; // @[TopModule.scala 192:48]
  wire [32:0] ConstUnit3_io_outputs_0; // @[TopModule.scala 192:48]
  wire [31:0] ConstUnit4_io_cfg; // @[TopModule.scala 192:48]
  wire [32:0] ConstUnit4_io_outputs_0; // @[TopModule.scala 192:48]
  wire [31:0] ConstUnit5_io_cfg; // @[TopModule.scala 192:48]
  wire [32:0] ConstUnit5_io_outputs_0; // @[TopModule.scala 192:48]
  wire [31:0] ConstUnit6_io_cfg; // @[TopModule.scala 192:48]
  wire [32:0] ConstUnit6_io_outputs_0; // @[TopModule.scala 192:48]
  wire [31:0] ConstUnit7_io_cfg; // @[TopModule.scala 192:48]
  wire [32:0] ConstUnit7_io_outputs_0; // @[TopModule.scala 192:48]
  wire [4:0] MUX0_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_18; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_19; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_20; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_21; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_22; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_23; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX1_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_18; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_19; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_20; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_21; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_22; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_23; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX2_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_18; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_19; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_20; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_21; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_22; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_23; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX3_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_18; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_19; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_20; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_21; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_22; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_23; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX4_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_18; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_19; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_20; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_21; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_22; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_23; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX5_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_18; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_19; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_20; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_21; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_22; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_23; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX6_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_18; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_19; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_20; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_21; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_22; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_23; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX7_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_18; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_19; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_20; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_21; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_22; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_23; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX8_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_18; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_19; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_20; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_21; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_22; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_23; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_24; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX9_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_18; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_19; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_20; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_21; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_22; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_23; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_24; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX10_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_18; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_19; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_20; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_21; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_22; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_23; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_24; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX11_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_18; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_19; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_20; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_21; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_22; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_23; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_24; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX12_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_18; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_19; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_20; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_21; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_22; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_23; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_24; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX13_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_18; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_19; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_20; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_21; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_22; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_23; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_24; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX14_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_18; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_19; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_20; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_21; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_22; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_23; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_24; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_outputs_0; // @[TopModule.scala 199:48]
  wire [4:0] MUX15_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_9; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_10; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_11; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_12; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_13; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_14; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_15; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_16; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_17; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_18; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_19; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_20; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_21; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_22; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_23; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_24; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_outputs_0; // @[TopModule.scala 199:48]
  wire  MUXR0_clock; // @[TopModule.scala 205:48]
  wire  MUXR0_reset; // @[TopModule.scala 205:48]
  wire [4:0] MUXR0_io_cfg; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_0; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_1; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_2; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_3; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_4; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_5; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_6; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_7; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_8; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_9; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_10; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_11; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_12; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_13; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_14; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_15; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_16; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_17; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_18; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_19; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_20; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_21; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_22; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_inputs_23; // @[TopModule.scala 205:48]
  wire [32:0] MUXR0_io_outputs_0; // @[TopModule.scala 205:48]
  wire  CfgMem_clock; // @[TopModule.scala 232:29]
  wire  CfgMem_reset; // @[TopModule.scala 232:29]
  wire  CfgMem_io_cfgEn; // @[TopModule.scala 232:29]
  wire [3:0] CfgMem_io_cfgAddr; // @[TopModule.scala 232:29]
  wire [31:0] CfgMem_io_cfgData; // @[TopModule.scala 232:29]
  wire [340:0] CfgMem_io_cfgOut; // @[TopModule.scala 232:29]
  ConstUnit0 ConstUnit0 ( // @[TopModule.scala 192:48]
    .io_cfg(ConstUnit0_io_cfg),
    .io_outputs_0(ConstUnit0_io_outputs_0)
  );
  ConstUnit0 ConstUnit1 ( // @[TopModule.scala 192:48]
    .io_cfg(ConstUnit1_io_cfg),
    .io_outputs_0(ConstUnit1_io_outputs_0)
  );
  ConstUnit0 ConstUnit2 ( // @[TopModule.scala 192:48]
    .io_cfg(ConstUnit2_io_cfg),
    .io_outputs_0(ConstUnit2_io_outputs_0)
  );
  ConstUnit0 ConstUnit3 ( // @[TopModule.scala 192:48]
    .io_cfg(ConstUnit3_io_cfg),
    .io_outputs_0(ConstUnit3_io_outputs_0)
  );
  ConstUnit0 ConstUnit4 ( // @[TopModule.scala 192:48]
    .io_cfg(ConstUnit4_io_cfg),
    .io_outputs_0(ConstUnit4_io_outputs_0)
  );
  ConstUnit0 ConstUnit5 ( // @[TopModule.scala 192:48]
    .io_cfg(ConstUnit5_io_cfg),
    .io_outputs_0(ConstUnit5_io_outputs_0)
  );
  ConstUnit0 ConstUnit6 ( // @[TopModule.scala 192:48]
    .io_cfg(ConstUnit6_io_cfg),
    .io_outputs_0(ConstUnit6_io_outputs_0)
  );
  ConstUnit0 ConstUnit7 ( // @[TopModule.scala 192:48]
    .io_cfg(ConstUnit7_io_cfg),
    .io_outputs_0(ConstUnit7_io_outputs_0)
  );
  MUX0_1 MUX0 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX0_io_cfg),
    .io_inputs_0(MUX0_io_inputs_0),
    .io_inputs_1(MUX0_io_inputs_1),
    .io_inputs_2(MUX0_io_inputs_2),
    .io_inputs_3(MUX0_io_inputs_3),
    .io_inputs_4(MUX0_io_inputs_4),
    .io_inputs_5(MUX0_io_inputs_5),
    .io_inputs_6(MUX0_io_inputs_6),
    .io_inputs_7(MUX0_io_inputs_7),
    .io_inputs_8(MUX0_io_inputs_8),
    .io_inputs_9(MUX0_io_inputs_9),
    .io_inputs_10(MUX0_io_inputs_10),
    .io_inputs_11(MUX0_io_inputs_11),
    .io_inputs_12(MUX0_io_inputs_12),
    .io_inputs_13(MUX0_io_inputs_13),
    .io_inputs_14(MUX0_io_inputs_14),
    .io_inputs_15(MUX0_io_inputs_15),
    .io_inputs_16(MUX0_io_inputs_16),
    .io_inputs_17(MUX0_io_inputs_17),
    .io_inputs_18(MUX0_io_inputs_18),
    .io_inputs_19(MUX0_io_inputs_19),
    .io_inputs_20(MUX0_io_inputs_20),
    .io_inputs_21(MUX0_io_inputs_21),
    .io_inputs_22(MUX0_io_inputs_22),
    .io_inputs_23(MUX0_io_inputs_23),
    .io_outputs_0(MUX0_io_outputs_0)
  );
  MUX0_1 MUX1 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX1_io_cfg),
    .io_inputs_0(MUX1_io_inputs_0),
    .io_inputs_1(MUX1_io_inputs_1),
    .io_inputs_2(MUX1_io_inputs_2),
    .io_inputs_3(MUX1_io_inputs_3),
    .io_inputs_4(MUX1_io_inputs_4),
    .io_inputs_5(MUX1_io_inputs_5),
    .io_inputs_6(MUX1_io_inputs_6),
    .io_inputs_7(MUX1_io_inputs_7),
    .io_inputs_8(MUX1_io_inputs_8),
    .io_inputs_9(MUX1_io_inputs_9),
    .io_inputs_10(MUX1_io_inputs_10),
    .io_inputs_11(MUX1_io_inputs_11),
    .io_inputs_12(MUX1_io_inputs_12),
    .io_inputs_13(MUX1_io_inputs_13),
    .io_inputs_14(MUX1_io_inputs_14),
    .io_inputs_15(MUX1_io_inputs_15),
    .io_inputs_16(MUX1_io_inputs_16),
    .io_inputs_17(MUX1_io_inputs_17),
    .io_inputs_18(MUX1_io_inputs_18),
    .io_inputs_19(MUX1_io_inputs_19),
    .io_inputs_20(MUX1_io_inputs_20),
    .io_inputs_21(MUX1_io_inputs_21),
    .io_inputs_22(MUX1_io_inputs_22),
    .io_inputs_23(MUX1_io_inputs_23),
    .io_outputs_0(MUX1_io_outputs_0)
  );
  MUX0_1 MUX2 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX2_io_cfg),
    .io_inputs_0(MUX2_io_inputs_0),
    .io_inputs_1(MUX2_io_inputs_1),
    .io_inputs_2(MUX2_io_inputs_2),
    .io_inputs_3(MUX2_io_inputs_3),
    .io_inputs_4(MUX2_io_inputs_4),
    .io_inputs_5(MUX2_io_inputs_5),
    .io_inputs_6(MUX2_io_inputs_6),
    .io_inputs_7(MUX2_io_inputs_7),
    .io_inputs_8(MUX2_io_inputs_8),
    .io_inputs_9(MUX2_io_inputs_9),
    .io_inputs_10(MUX2_io_inputs_10),
    .io_inputs_11(MUX2_io_inputs_11),
    .io_inputs_12(MUX2_io_inputs_12),
    .io_inputs_13(MUX2_io_inputs_13),
    .io_inputs_14(MUX2_io_inputs_14),
    .io_inputs_15(MUX2_io_inputs_15),
    .io_inputs_16(MUX2_io_inputs_16),
    .io_inputs_17(MUX2_io_inputs_17),
    .io_inputs_18(MUX2_io_inputs_18),
    .io_inputs_19(MUX2_io_inputs_19),
    .io_inputs_20(MUX2_io_inputs_20),
    .io_inputs_21(MUX2_io_inputs_21),
    .io_inputs_22(MUX2_io_inputs_22),
    .io_inputs_23(MUX2_io_inputs_23),
    .io_outputs_0(MUX2_io_outputs_0)
  );
  MUX0_1 MUX3 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX3_io_cfg),
    .io_inputs_0(MUX3_io_inputs_0),
    .io_inputs_1(MUX3_io_inputs_1),
    .io_inputs_2(MUX3_io_inputs_2),
    .io_inputs_3(MUX3_io_inputs_3),
    .io_inputs_4(MUX3_io_inputs_4),
    .io_inputs_5(MUX3_io_inputs_5),
    .io_inputs_6(MUX3_io_inputs_6),
    .io_inputs_7(MUX3_io_inputs_7),
    .io_inputs_8(MUX3_io_inputs_8),
    .io_inputs_9(MUX3_io_inputs_9),
    .io_inputs_10(MUX3_io_inputs_10),
    .io_inputs_11(MUX3_io_inputs_11),
    .io_inputs_12(MUX3_io_inputs_12),
    .io_inputs_13(MUX3_io_inputs_13),
    .io_inputs_14(MUX3_io_inputs_14),
    .io_inputs_15(MUX3_io_inputs_15),
    .io_inputs_16(MUX3_io_inputs_16),
    .io_inputs_17(MUX3_io_inputs_17),
    .io_inputs_18(MUX3_io_inputs_18),
    .io_inputs_19(MUX3_io_inputs_19),
    .io_inputs_20(MUX3_io_inputs_20),
    .io_inputs_21(MUX3_io_inputs_21),
    .io_inputs_22(MUX3_io_inputs_22),
    .io_inputs_23(MUX3_io_inputs_23),
    .io_outputs_0(MUX3_io_outputs_0)
  );
  MUX0_1 MUX4 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX4_io_cfg),
    .io_inputs_0(MUX4_io_inputs_0),
    .io_inputs_1(MUX4_io_inputs_1),
    .io_inputs_2(MUX4_io_inputs_2),
    .io_inputs_3(MUX4_io_inputs_3),
    .io_inputs_4(MUX4_io_inputs_4),
    .io_inputs_5(MUX4_io_inputs_5),
    .io_inputs_6(MUX4_io_inputs_6),
    .io_inputs_7(MUX4_io_inputs_7),
    .io_inputs_8(MUX4_io_inputs_8),
    .io_inputs_9(MUX4_io_inputs_9),
    .io_inputs_10(MUX4_io_inputs_10),
    .io_inputs_11(MUX4_io_inputs_11),
    .io_inputs_12(MUX4_io_inputs_12),
    .io_inputs_13(MUX4_io_inputs_13),
    .io_inputs_14(MUX4_io_inputs_14),
    .io_inputs_15(MUX4_io_inputs_15),
    .io_inputs_16(MUX4_io_inputs_16),
    .io_inputs_17(MUX4_io_inputs_17),
    .io_inputs_18(MUX4_io_inputs_18),
    .io_inputs_19(MUX4_io_inputs_19),
    .io_inputs_20(MUX4_io_inputs_20),
    .io_inputs_21(MUX4_io_inputs_21),
    .io_inputs_22(MUX4_io_inputs_22),
    .io_inputs_23(MUX4_io_inputs_23),
    .io_outputs_0(MUX4_io_outputs_0)
  );
  MUX0_1 MUX5 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX5_io_cfg),
    .io_inputs_0(MUX5_io_inputs_0),
    .io_inputs_1(MUX5_io_inputs_1),
    .io_inputs_2(MUX5_io_inputs_2),
    .io_inputs_3(MUX5_io_inputs_3),
    .io_inputs_4(MUX5_io_inputs_4),
    .io_inputs_5(MUX5_io_inputs_5),
    .io_inputs_6(MUX5_io_inputs_6),
    .io_inputs_7(MUX5_io_inputs_7),
    .io_inputs_8(MUX5_io_inputs_8),
    .io_inputs_9(MUX5_io_inputs_9),
    .io_inputs_10(MUX5_io_inputs_10),
    .io_inputs_11(MUX5_io_inputs_11),
    .io_inputs_12(MUX5_io_inputs_12),
    .io_inputs_13(MUX5_io_inputs_13),
    .io_inputs_14(MUX5_io_inputs_14),
    .io_inputs_15(MUX5_io_inputs_15),
    .io_inputs_16(MUX5_io_inputs_16),
    .io_inputs_17(MUX5_io_inputs_17),
    .io_inputs_18(MUX5_io_inputs_18),
    .io_inputs_19(MUX5_io_inputs_19),
    .io_inputs_20(MUX5_io_inputs_20),
    .io_inputs_21(MUX5_io_inputs_21),
    .io_inputs_22(MUX5_io_inputs_22),
    .io_inputs_23(MUX5_io_inputs_23),
    .io_outputs_0(MUX5_io_outputs_0)
  );
  MUX0_1 MUX6 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX6_io_cfg),
    .io_inputs_0(MUX6_io_inputs_0),
    .io_inputs_1(MUX6_io_inputs_1),
    .io_inputs_2(MUX6_io_inputs_2),
    .io_inputs_3(MUX6_io_inputs_3),
    .io_inputs_4(MUX6_io_inputs_4),
    .io_inputs_5(MUX6_io_inputs_5),
    .io_inputs_6(MUX6_io_inputs_6),
    .io_inputs_7(MUX6_io_inputs_7),
    .io_inputs_8(MUX6_io_inputs_8),
    .io_inputs_9(MUX6_io_inputs_9),
    .io_inputs_10(MUX6_io_inputs_10),
    .io_inputs_11(MUX6_io_inputs_11),
    .io_inputs_12(MUX6_io_inputs_12),
    .io_inputs_13(MUX6_io_inputs_13),
    .io_inputs_14(MUX6_io_inputs_14),
    .io_inputs_15(MUX6_io_inputs_15),
    .io_inputs_16(MUX6_io_inputs_16),
    .io_inputs_17(MUX6_io_inputs_17),
    .io_inputs_18(MUX6_io_inputs_18),
    .io_inputs_19(MUX6_io_inputs_19),
    .io_inputs_20(MUX6_io_inputs_20),
    .io_inputs_21(MUX6_io_inputs_21),
    .io_inputs_22(MUX6_io_inputs_22),
    .io_inputs_23(MUX6_io_inputs_23),
    .io_outputs_0(MUX6_io_outputs_0)
  );
  MUX0_1 MUX7 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX7_io_cfg),
    .io_inputs_0(MUX7_io_inputs_0),
    .io_inputs_1(MUX7_io_inputs_1),
    .io_inputs_2(MUX7_io_inputs_2),
    .io_inputs_3(MUX7_io_inputs_3),
    .io_inputs_4(MUX7_io_inputs_4),
    .io_inputs_5(MUX7_io_inputs_5),
    .io_inputs_6(MUX7_io_inputs_6),
    .io_inputs_7(MUX7_io_inputs_7),
    .io_inputs_8(MUX7_io_inputs_8),
    .io_inputs_9(MUX7_io_inputs_9),
    .io_inputs_10(MUX7_io_inputs_10),
    .io_inputs_11(MUX7_io_inputs_11),
    .io_inputs_12(MUX7_io_inputs_12),
    .io_inputs_13(MUX7_io_inputs_13),
    .io_inputs_14(MUX7_io_inputs_14),
    .io_inputs_15(MUX7_io_inputs_15),
    .io_inputs_16(MUX7_io_inputs_16),
    .io_inputs_17(MUX7_io_inputs_17),
    .io_inputs_18(MUX7_io_inputs_18),
    .io_inputs_19(MUX7_io_inputs_19),
    .io_inputs_20(MUX7_io_inputs_20),
    .io_inputs_21(MUX7_io_inputs_21),
    .io_inputs_22(MUX7_io_inputs_22),
    .io_inputs_23(MUX7_io_inputs_23),
    .io_outputs_0(MUX7_io_outputs_0)
  );
  MUX8_1 MUX8 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX8_io_cfg),
    .io_inputs_0(MUX8_io_inputs_0),
    .io_inputs_1(MUX8_io_inputs_1),
    .io_inputs_2(MUX8_io_inputs_2),
    .io_inputs_3(MUX8_io_inputs_3),
    .io_inputs_4(MUX8_io_inputs_4),
    .io_inputs_5(MUX8_io_inputs_5),
    .io_inputs_6(MUX8_io_inputs_6),
    .io_inputs_7(MUX8_io_inputs_7),
    .io_inputs_8(MUX8_io_inputs_8),
    .io_inputs_9(MUX8_io_inputs_9),
    .io_inputs_10(MUX8_io_inputs_10),
    .io_inputs_11(MUX8_io_inputs_11),
    .io_inputs_12(MUX8_io_inputs_12),
    .io_inputs_13(MUX8_io_inputs_13),
    .io_inputs_14(MUX8_io_inputs_14),
    .io_inputs_15(MUX8_io_inputs_15),
    .io_inputs_16(MUX8_io_inputs_16),
    .io_inputs_17(MUX8_io_inputs_17),
    .io_inputs_18(MUX8_io_inputs_18),
    .io_inputs_19(MUX8_io_inputs_19),
    .io_inputs_20(MUX8_io_inputs_20),
    .io_inputs_21(MUX8_io_inputs_21),
    .io_inputs_22(MUX8_io_inputs_22),
    .io_inputs_23(MUX8_io_inputs_23),
    .io_inputs_24(MUX8_io_inputs_24),
    .io_outputs_0(MUX8_io_outputs_0)
  );
  MUX8_1 MUX9 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX9_io_cfg),
    .io_inputs_0(MUX9_io_inputs_0),
    .io_inputs_1(MUX9_io_inputs_1),
    .io_inputs_2(MUX9_io_inputs_2),
    .io_inputs_3(MUX9_io_inputs_3),
    .io_inputs_4(MUX9_io_inputs_4),
    .io_inputs_5(MUX9_io_inputs_5),
    .io_inputs_6(MUX9_io_inputs_6),
    .io_inputs_7(MUX9_io_inputs_7),
    .io_inputs_8(MUX9_io_inputs_8),
    .io_inputs_9(MUX9_io_inputs_9),
    .io_inputs_10(MUX9_io_inputs_10),
    .io_inputs_11(MUX9_io_inputs_11),
    .io_inputs_12(MUX9_io_inputs_12),
    .io_inputs_13(MUX9_io_inputs_13),
    .io_inputs_14(MUX9_io_inputs_14),
    .io_inputs_15(MUX9_io_inputs_15),
    .io_inputs_16(MUX9_io_inputs_16),
    .io_inputs_17(MUX9_io_inputs_17),
    .io_inputs_18(MUX9_io_inputs_18),
    .io_inputs_19(MUX9_io_inputs_19),
    .io_inputs_20(MUX9_io_inputs_20),
    .io_inputs_21(MUX9_io_inputs_21),
    .io_inputs_22(MUX9_io_inputs_22),
    .io_inputs_23(MUX9_io_inputs_23),
    .io_inputs_24(MUX9_io_inputs_24),
    .io_outputs_0(MUX9_io_outputs_0)
  );
  MUX8_1 MUX10 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX10_io_cfg),
    .io_inputs_0(MUX10_io_inputs_0),
    .io_inputs_1(MUX10_io_inputs_1),
    .io_inputs_2(MUX10_io_inputs_2),
    .io_inputs_3(MUX10_io_inputs_3),
    .io_inputs_4(MUX10_io_inputs_4),
    .io_inputs_5(MUX10_io_inputs_5),
    .io_inputs_6(MUX10_io_inputs_6),
    .io_inputs_7(MUX10_io_inputs_7),
    .io_inputs_8(MUX10_io_inputs_8),
    .io_inputs_9(MUX10_io_inputs_9),
    .io_inputs_10(MUX10_io_inputs_10),
    .io_inputs_11(MUX10_io_inputs_11),
    .io_inputs_12(MUX10_io_inputs_12),
    .io_inputs_13(MUX10_io_inputs_13),
    .io_inputs_14(MUX10_io_inputs_14),
    .io_inputs_15(MUX10_io_inputs_15),
    .io_inputs_16(MUX10_io_inputs_16),
    .io_inputs_17(MUX10_io_inputs_17),
    .io_inputs_18(MUX10_io_inputs_18),
    .io_inputs_19(MUX10_io_inputs_19),
    .io_inputs_20(MUX10_io_inputs_20),
    .io_inputs_21(MUX10_io_inputs_21),
    .io_inputs_22(MUX10_io_inputs_22),
    .io_inputs_23(MUX10_io_inputs_23),
    .io_inputs_24(MUX10_io_inputs_24),
    .io_outputs_0(MUX10_io_outputs_0)
  );
  MUX8_1 MUX11 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX11_io_cfg),
    .io_inputs_0(MUX11_io_inputs_0),
    .io_inputs_1(MUX11_io_inputs_1),
    .io_inputs_2(MUX11_io_inputs_2),
    .io_inputs_3(MUX11_io_inputs_3),
    .io_inputs_4(MUX11_io_inputs_4),
    .io_inputs_5(MUX11_io_inputs_5),
    .io_inputs_6(MUX11_io_inputs_6),
    .io_inputs_7(MUX11_io_inputs_7),
    .io_inputs_8(MUX11_io_inputs_8),
    .io_inputs_9(MUX11_io_inputs_9),
    .io_inputs_10(MUX11_io_inputs_10),
    .io_inputs_11(MUX11_io_inputs_11),
    .io_inputs_12(MUX11_io_inputs_12),
    .io_inputs_13(MUX11_io_inputs_13),
    .io_inputs_14(MUX11_io_inputs_14),
    .io_inputs_15(MUX11_io_inputs_15),
    .io_inputs_16(MUX11_io_inputs_16),
    .io_inputs_17(MUX11_io_inputs_17),
    .io_inputs_18(MUX11_io_inputs_18),
    .io_inputs_19(MUX11_io_inputs_19),
    .io_inputs_20(MUX11_io_inputs_20),
    .io_inputs_21(MUX11_io_inputs_21),
    .io_inputs_22(MUX11_io_inputs_22),
    .io_inputs_23(MUX11_io_inputs_23),
    .io_inputs_24(MUX11_io_inputs_24),
    .io_outputs_0(MUX11_io_outputs_0)
  );
  MUX8_1 MUX12 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX12_io_cfg),
    .io_inputs_0(MUX12_io_inputs_0),
    .io_inputs_1(MUX12_io_inputs_1),
    .io_inputs_2(MUX12_io_inputs_2),
    .io_inputs_3(MUX12_io_inputs_3),
    .io_inputs_4(MUX12_io_inputs_4),
    .io_inputs_5(MUX12_io_inputs_5),
    .io_inputs_6(MUX12_io_inputs_6),
    .io_inputs_7(MUX12_io_inputs_7),
    .io_inputs_8(MUX12_io_inputs_8),
    .io_inputs_9(MUX12_io_inputs_9),
    .io_inputs_10(MUX12_io_inputs_10),
    .io_inputs_11(MUX12_io_inputs_11),
    .io_inputs_12(MUX12_io_inputs_12),
    .io_inputs_13(MUX12_io_inputs_13),
    .io_inputs_14(MUX12_io_inputs_14),
    .io_inputs_15(MUX12_io_inputs_15),
    .io_inputs_16(MUX12_io_inputs_16),
    .io_inputs_17(MUX12_io_inputs_17),
    .io_inputs_18(MUX12_io_inputs_18),
    .io_inputs_19(MUX12_io_inputs_19),
    .io_inputs_20(MUX12_io_inputs_20),
    .io_inputs_21(MUX12_io_inputs_21),
    .io_inputs_22(MUX12_io_inputs_22),
    .io_inputs_23(MUX12_io_inputs_23),
    .io_inputs_24(MUX12_io_inputs_24),
    .io_outputs_0(MUX12_io_outputs_0)
  );
  MUX8_1 MUX13 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX13_io_cfg),
    .io_inputs_0(MUX13_io_inputs_0),
    .io_inputs_1(MUX13_io_inputs_1),
    .io_inputs_2(MUX13_io_inputs_2),
    .io_inputs_3(MUX13_io_inputs_3),
    .io_inputs_4(MUX13_io_inputs_4),
    .io_inputs_5(MUX13_io_inputs_5),
    .io_inputs_6(MUX13_io_inputs_6),
    .io_inputs_7(MUX13_io_inputs_7),
    .io_inputs_8(MUX13_io_inputs_8),
    .io_inputs_9(MUX13_io_inputs_9),
    .io_inputs_10(MUX13_io_inputs_10),
    .io_inputs_11(MUX13_io_inputs_11),
    .io_inputs_12(MUX13_io_inputs_12),
    .io_inputs_13(MUX13_io_inputs_13),
    .io_inputs_14(MUX13_io_inputs_14),
    .io_inputs_15(MUX13_io_inputs_15),
    .io_inputs_16(MUX13_io_inputs_16),
    .io_inputs_17(MUX13_io_inputs_17),
    .io_inputs_18(MUX13_io_inputs_18),
    .io_inputs_19(MUX13_io_inputs_19),
    .io_inputs_20(MUX13_io_inputs_20),
    .io_inputs_21(MUX13_io_inputs_21),
    .io_inputs_22(MUX13_io_inputs_22),
    .io_inputs_23(MUX13_io_inputs_23),
    .io_inputs_24(MUX13_io_inputs_24),
    .io_outputs_0(MUX13_io_outputs_0)
  );
  MUX8_1 MUX14 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX14_io_cfg),
    .io_inputs_0(MUX14_io_inputs_0),
    .io_inputs_1(MUX14_io_inputs_1),
    .io_inputs_2(MUX14_io_inputs_2),
    .io_inputs_3(MUX14_io_inputs_3),
    .io_inputs_4(MUX14_io_inputs_4),
    .io_inputs_5(MUX14_io_inputs_5),
    .io_inputs_6(MUX14_io_inputs_6),
    .io_inputs_7(MUX14_io_inputs_7),
    .io_inputs_8(MUX14_io_inputs_8),
    .io_inputs_9(MUX14_io_inputs_9),
    .io_inputs_10(MUX14_io_inputs_10),
    .io_inputs_11(MUX14_io_inputs_11),
    .io_inputs_12(MUX14_io_inputs_12),
    .io_inputs_13(MUX14_io_inputs_13),
    .io_inputs_14(MUX14_io_inputs_14),
    .io_inputs_15(MUX14_io_inputs_15),
    .io_inputs_16(MUX14_io_inputs_16),
    .io_inputs_17(MUX14_io_inputs_17),
    .io_inputs_18(MUX14_io_inputs_18),
    .io_inputs_19(MUX14_io_inputs_19),
    .io_inputs_20(MUX14_io_inputs_20),
    .io_inputs_21(MUX14_io_inputs_21),
    .io_inputs_22(MUX14_io_inputs_22),
    .io_inputs_23(MUX14_io_inputs_23),
    .io_inputs_24(MUX14_io_inputs_24),
    .io_outputs_0(MUX14_io_outputs_0)
  );
  MUX8_1 MUX15 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX15_io_cfg),
    .io_inputs_0(MUX15_io_inputs_0),
    .io_inputs_1(MUX15_io_inputs_1),
    .io_inputs_2(MUX15_io_inputs_2),
    .io_inputs_3(MUX15_io_inputs_3),
    .io_inputs_4(MUX15_io_inputs_4),
    .io_inputs_5(MUX15_io_inputs_5),
    .io_inputs_6(MUX15_io_inputs_6),
    .io_inputs_7(MUX15_io_inputs_7),
    .io_inputs_8(MUX15_io_inputs_8),
    .io_inputs_9(MUX15_io_inputs_9),
    .io_inputs_10(MUX15_io_inputs_10),
    .io_inputs_11(MUX15_io_inputs_11),
    .io_inputs_12(MUX15_io_inputs_12),
    .io_inputs_13(MUX15_io_inputs_13),
    .io_inputs_14(MUX15_io_inputs_14),
    .io_inputs_15(MUX15_io_inputs_15),
    .io_inputs_16(MUX15_io_inputs_16),
    .io_inputs_17(MUX15_io_inputs_17),
    .io_inputs_18(MUX15_io_inputs_18),
    .io_inputs_19(MUX15_io_inputs_19),
    .io_inputs_20(MUX15_io_inputs_20),
    .io_inputs_21(MUX15_io_inputs_21),
    .io_inputs_22(MUX15_io_inputs_22),
    .io_inputs_23(MUX15_io_inputs_23),
    .io_inputs_24(MUX15_io_inputs_24),
    .io_outputs_0(MUX15_io_outputs_0)
  );
  MUXR0_1 MUXR0 ( // @[TopModule.scala 205:48]
    .clock(MUXR0_clock),
    .reset(MUXR0_reset),
    .io_cfg(MUXR0_io_cfg),
    .io_inputs_0(MUXR0_io_inputs_0),
    .io_inputs_1(MUXR0_io_inputs_1),
    .io_inputs_2(MUXR0_io_inputs_2),
    .io_inputs_3(MUXR0_io_inputs_3),
    .io_inputs_4(MUXR0_io_inputs_4),
    .io_inputs_5(MUXR0_io_inputs_5),
    .io_inputs_6(MUXR0_io_inputs_6),
    .io_inputs_7(MUXR0_io_inputs_7),
    .io_inputs_8(MUXR0_io_inputs_8),
    .io_inputs_9(MUXR0_io_inputs_9),
    .io_inputs_10(MUXR0_io_inputs_10),
    .io_inputs_11(MUXR0_io_inputs_11),
    .io_inputs_12(MUXR0_io_inputs_12),
    .io_inputs_13(MUXR0_io_inputs_13),
    .io_inputs_14(MUXR0_io_inputs_14),
    .io_inputs_15(MUXR0_io_inputs_15),
    .io_inputs_16(MUXR0_io_inputs_16),
    .io_inputs_17(MUXR0_io_inputs_17),
    .io_inputs_18(MUXR0_io_inputs_18),
    .io_inputs_19(MUXR0_io_inputs_19),
    .io_inputs_20(MUXR0_io_inputs_20),
    .io_inputs_21(MUXR0_io_inputs_21),
    .io_inputs_22(MUXR0_io_inputs_22),
    .io_inputs_23(MUXR0_io_inputs_23),
    .io_outputs_0(MUXR0_io_outputs_0)
  );
  CfgMem_16 CfgMem ( // @[TopModule.scala 232:29]
    .clock(CfgMem_clock),
    .reset(CfgMem_reset),
    .io_cfgEn(CfgMem_io_cfgEn),
    .io_cfgAddr(CfgMem_io_cfgAddr),
    .io_cfgData(CfgMem_io_cfgData),
    .io_cfgOut(CfgMem_io_cfgOut)
  );
  assign io_outputs_0 = MUXR0_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_1 = MUX0_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_2 = MUX1_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_3 = MUX2_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_4 = MUX3_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_5 = MUX4_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_6 = MUX5_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_7 = MUX6_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_8 = MUX7_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_9 = MUX8_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_10 = MUX9_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_11 = MUX10_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_12 = MUX11_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_13 = MUX12_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_14 = MUX13_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_15 = MUX14_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_16 = MUX15_io_outputs_0; // @[TopModule.scala 392:22]
  assign ConstUnit0_io_cfg = CfgMem_io_cfgOut[31:0]; // @[TopModule.scala 259:94]
  assign ConstUnit1_io_cfg = CfgMem_io_cfgOut[63:32]; // @[TopModule.scala 259:94]
  assign ConstUnit2_io_cfg = CfgMem_io_cfgOut[95:64]; // @[TopModule.scala 259:94]
  assign ConstUnit3_io_cfg = CfgMem_io_cfgOut[127:96]; // @[TopModule.scala 259:94]
  assign ConstUnit4_io_cfg = CfgMem_io_cfgOut[159:128]; // @[TopModule.scala 259:94]
  assign ConstUnit5_io_cfg = CfgMem_io_cfgOut[191:160]; // @[TopModule.scala 259:94]
  assign ConstUnit6_io_cfg = CfgMem_io_cfgOut[223:192]; // @[TopModule.scala 259:94]
  assign ConstUnit7_io_cfg = CfgMem_io_cfgOut[255:224]; // @[TopModule.scala 259:94]
  assign MUX0_io_cfg = CfgMem_io_cfgOut[260:256]; // @[TopModule.scala 261:98]
  assign MUX0_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_17 = io_inputs_17; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_18 = io_inputs_18; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_19 = io_inputs_19; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_20 = io_inputs_20; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_21 = io_inputs_21; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_22 = io_inputs_22; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_23 = io_inputs_23; // @[TopModule.scala 392:22]
  assign MUX1_io_cfg = CfgMem_io_cfgOut[265:261]; // @[TopModule.scala 261:98]
  assign MUX1_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_17 = io_inputs_17; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_18 = io_inputs_18; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_19 = io_inputs_19; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_20 = io_inputs_20; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_21 = io_inputs_21; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_22 = io_inputs_22; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_23 = io_inputs_23; // @[TopModule.scala 392:22]
  assign MUX2_io_cfg = CfgMem_io_cfgOut[270:266]; // @[TopModule.scala 261:98]
  assign MUX2_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_17 = io_inputs_17; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_18 = io_inputs_18; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_19 = io_inputs_19; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_20 = io_inputs_20; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_21 = io_inputs_21; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_22 = io_inputs_22; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_23 = io_inputs_23; // @[TopModule.scala 392:22]
  assign MUX3_io_cfg = CfgMem_io_cfgOut[275:271]; // @[TopModule.scala 261:98]
  assign MUX3_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_17 = io_inputs_17; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_18 = io_inputs_18; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_19 = io_inputs_19; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_20 = io_inputs_20; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_21 = io_inputs_21; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_22 = io_inputs_22; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_23 = io_inputs_23; // @[TopModule.scala 392:22]
  assign MUX4_io_cfg = CfgMem_io_cfgOut[280:276]; // @[TopModule.scala 261:98]
  assign MUX4_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_17 = io_inputs_17; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_18 = io_inputs_18; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_19 = io_inputs_19; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_20 = io_inputs_20; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_21 = io_inputs_21; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_22 = io_inputs_22; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_23 = io_inputs_23; // @[TopModule.scala 392:22]
  assign MUX5_io_cfg = CfgMem_io_cfgOut[285:281]; // @[TopModule.scala 261:98]
  assign MUX5_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_17 = io_inputs_17; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_18 = io_inputs_18; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_19 = io_inputs_19; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_20 = io_inputs_20; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_21 = io_inputs_21; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_22 = io_inputs_22; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_23 = io_inputs_23; // @[TopModule.scala 392:22]
  assign MUX6_io_cfg = CfgMem_io_cfgOut[290:286]; // @[TopModule.scala 261:98]
  assign MUX6_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_17 = io_inputs_17; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_18 = io_inputs_18; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_19 = io_inputs_19; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_20 = io_inputs_20; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_21 = io_inputs_21; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_22 = io_inputs_22; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_23 = io_inputs_23; // @[TopModule.scala 392:22]
  assign MUX7_io_cfg = CfgMem_io_cfgOut[295:291]; // @[TopModule.scala 261:98]
  assign MUX7_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_17 = io_inputs_17; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_18 = io_inputs_18; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_19 = io_inputs_19; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_20 = io_inputs_20; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_21 = io_inputs_21; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_22 = io_inputs_22; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_23 = io_inputs_23; // @[TopModule.scala 392:22]
  assign MUX8_io_cfg = CfgMem_io_cfgOut[300:296]; // @[TopModule.scala 261:98]
  assign MUX8_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_17 = io_inputs_17; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_18 = io_inputs_18; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_19 = io_inputs_19; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_20 = io_inputs_20; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_21 = io_inputs_21; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_22 = io_inputs_22; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_23 = io_inputs_23; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_24 = ConstUnit0_io_outputs_0; // @[TopModule.scala 392:22]
  assign MUX9_io_cfg = CfgMem_io_cfgOut[305:301]; // @[TopModule.scala 261:98]
  assign MUX9_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_17 = io_inputs_17; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_18 = io_inputs_18; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_19 = io_inputs_19; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_20 = io_inputs_20; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_21 = io_inputs_21; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_22 = io_inputs_22; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_23 = io_inputs_23; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_24 = ConstUnit1_io_outputs_0; // @[TopModule.scala 392:22]
  assign MUX10_io_cfg = CfgMem_io_cfgOut[310:306]; // @[TopModule.scala 261:98]
  assign MUX10_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_17 = io_inputs_17; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_18 = io_inputs_18; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_19 = io_inputs_19; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_20 = io_inputs_20; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_21 = io_inputs_21; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_22 = io_inputs_22; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_23 = io_inputs_23; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_24 = ConstUnit2_io_outputs_0; // @[TopModule.scala 392:22]
  assign MUX11_io_cfg = CfgMem_io_cfgOut[315:311]; // @[TopModule.scala 261:98]
  assign MUX11_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_17 = io_inputs_17; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_18 = io_inputs_18; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_19 = io_inputs_19; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_20 = io_inputs_20; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_21 = io_inputs_21; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_22 = io_inputs_22; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_23 = io_inputs_23; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_24 = ConstUnit3_io_outputs_0; // @[TopModule.scala 392:22]
  assign MUX12_io_cfg = CfgMem_io_cfgOut[320:316]; // @[TopModule.scala 261:98]
  assign MUX12_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_17 = io_inputs_17; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_18 = io_inputs_18; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_19 = io_inputs_19; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_20 = io_inputs_20; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_21 = io_inputs_21; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_22 = io_inputs_22; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_23 = io_inputs_23; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_24 = ConstUnit4_io_outputs_0; // @[TopModule.scala 392:22]
  assign MUX13_io_cfg = CfgMem_io_cfgOut[325:321]; // @[TopModule.scala 261:98]
  assign MUX13_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_17 = io_inputs_17; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_18 = io_inputs_18; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_19 = io_inputs_19; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_20 = io_inputs_20; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_21 = io_inputs_21; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_22 = io_inputs_22; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_23 = io_inputs_23; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_24 = ConstUnit5_io_outputs_0; // @[TopModule.scala 392:22]
  assign MUX14_io_cfg = CfgMem_io_cfgOut[330:326]; // @[TopModule.scala 261:98]
  assign MUX14_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_17 = io_inputs_17; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_18 = io_inputs_18; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_19 = io_inputs_19; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_20 = io_inputs_20; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_21 = io_inputs_21; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_22 = io_inputs_22; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_23 = io_inputs_23; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_24 = ConstUnit6_io_outputs_0; // @[TopModule.scala 392:22]
  assign MUX15_io_cfg = CfgMem_io_cfgOut[335:331]; // @[TopModule.scala 261:98]
  assign MUX15_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_17 = io_inputs_17; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_18 = io_inputs_18; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_19 = io_inputs_19; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_20 = io_inputs_20; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_21 = io_inputs_21; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_22 = io_inputs_22; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_23 = io_inputs_23; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_24 = ConstUnit7_io_outputs_0; // @[TopModule.scala 392:22]
  assign MUXR0_clock = clock;
  assign MUXR0_reset = reset;
  assign MUXR0_io_cfg = CfgMem_io_cfgOut[340:336]; // @[TopModule.scala 262:100]
  assign MUXR0_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_9 = io_inputs_9; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_10 = io_inputs_10; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_11 = io_inputs_11; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_12 = io_inputs_12; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_13 = io_inputs_13; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_14 = io_inputs_14; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_15 = io_inputs_15; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_16 = io_inputs_16; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_17 = io_inputs_17; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_18 = io_inputs_18; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_19 = io_inputs_19; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_20 = io_inputs_20; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_21 = io_inputs_21; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_22 = io_inputs_22; // @[TopModule.scala 392:22]
  assign MUXR0_io_inputs_23 = io_inputs_23; // @[TopModule.scala 392:22]
  assign CfgMem_clock = clock;
  assign CfgMem_reset = reset;
  assign CfgMem_io_cfgEn = io_cfgEn; // @[TopModule.scala 239:34]
  assign CfgMem_io_cfgAddr = io_cfgAddr; // @[TopModule.scala 244:30]
  assign CfgMem_io_cfgData = io_cfgData; // @[TopModule.scala 248:28]
endmodule
module MUX0_2(
  input  [3:0]  io_cfg,
  input  [32:0] io_inputs_0,
  input  [32:0] io_inputs_1,
  input  [32:0] io_inputs_2,
  input  [32:0] io_inputs_3,
  input  [32:0] io_inputs_4,
  input  [32:0] io_inputs_5,
  input  [32:0] io_inputs_6,
  input  [32:0] io_inputs_7,
  input  [32:0] io_inputs_8,
  output [32:0] io_outputs_0
);
  wire  _T = 4'h0 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_1 = _T ? io_inputs_0 : 33'h0; // @[Mux.scala 80:57]
  wire  _T_2 = 4'h1 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_3 = _T_2 ? io_inputs_1 : _T_1; // @[Mux.scala 80:57]
  wire  _T_4 = 4'h2 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_5 = _T_4 ? io_inputs_2 : _T_3; // @[Mux.scala 80:57]
  wire  _T_6 = 4'h3 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_7 = _T_6 ? io_inputs_3 : _T_5; // @[Mux.scala 80:57]
  wire  _T_8 = 4'h4 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_9 = _T_8 ? io_inputs_4 : _T_7; // @[Mux.scala 80:57]
  wire  _T_10 = 4'h5 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_11 = _T_10 ? io_inputs_5 : _T_9; // @[Mux.scala 80:57]
  wire  _T_12 = 4'h6 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_13 = _T_12 ? io_inputs_6 : _T_11; // @[Mux.scala 80:57]
  wire  _T_14 = 4'h7 == io_cfg; // @[Mux.scala 80:60]
  wire [32:0] _T_15 = _T_14 ? io_inputs_7 : _T_13; // @[Mux.scala 80:57]
  wire  _T_16 = 4'h8 == io_cfg; // @[Mux.scala 80:60]
  assign io_outputs_0 = _T_16 ? io_inputs_8 : _T_15; // @[Multiplexer.scala 16:17]
endmodule
module CfgMem_18(
  input         clock,
  input         reset,
  input         io_cfgEn,
  input         io_cfgAddr,
  input  [31:0] io_cfgData,
  output [63:0] io_cfgOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _T = ~io_cfgAddr; // @[CfgMem.scala 20:71]
  wire  _T_1 = io_cfgEn & _T; // @[CfgMem.scala 20:57]
  reg [31:0] outWire_0; // @[Reg.scala 27:20]
  wire  _T_4 = io_cfgEn & io_cfgAddr; // @[CfgMem.scala 20:57]
  reg [31:0] outWire_1; // @[Reg.scala 27:20]
  assign io_cfgOut = {outWire_1,outWire_0}; // @[CfgMem.scala 22:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  outWire_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  outWire_1 = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      outWire_0 <= 32'h0;
    end else if (_T_1) begin
      outWire_0 <= io_cfgData;
    end
    if (reset) begin
      outWire_1 <= 32'h0;
    end else if (_T_4) begin
      outWire_1 <= io_cfgData;
    end
  end
endmodule
module matrixFCdevice2(
  input         clock,
  input         reset,
  input         io_cfgEn,
  input  [3:0]  io_cfgAddr,
  input  [31:0] io_cfgData,
  input  [32:0] io_inputs_0,
  input  [32:0] io_inputs_1,
  input  [32:0] io_inputs_2,
  input  [32:0] io_inputs_3,
  input  [32:0] io_inputs_4,
  input  [32:0] io_inputs_5,
  input  [32:0] io_inputs_6,
  input  [32:0] io_inputs_7,
  input  [32:0] io_inputs_8,
  output [32:0] io_outputs_0,
  output [32:0] io_outputs_1,
  output [32:0] io_outputs_2,
  output [32:0] io_outputs_3,
  output [32:0] io_outputs_4,
  output [32:0] io_outputs_5,
  output [32:0] io_outputs_6,
  output [32:0] io_outputs_7,
  output [32:0] io_outputs_8,
  output [32:0] io_outputs_9,
  output [32:0] io_outputs_10,
  output [32:0] io_outputs_11,
  output [32:0] io_outputs_12,
  output [32:0] io_outputs_13,
  output [32:0] io_outputs_14,
  output [32:0] io_outputs_15
);
  wire [3:0] MUX0_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX0_io_outputs_0; // @[TopModule.scala 199:48]
  wire [3:0] MUX1_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX1_io_outputs_0; // @[TopModule.scala 199:48]
  wire [3:0] MUX2_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX2_io_outputs_0; // @[TopModule.scala 199:48]
  wire [3:0] MUX3_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX3_io_outputs_0; // @[TopModule.scala 199:48]
  wire [3:0] MUX4_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX4_io_outputs_0; // @[TopModule.scala 199:48]
  wire [3:0] MUX5_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX5_io_outputs_0; // @[TopModule.scala 199:48]
  wire [3:0] MUX6_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX6_io_outputs_0; // @[TopModule.scala 199:48]
  wire [3:0] MUX7_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX7_io_outputs_0; // @[TopModule.scala 199:48]
  wire [3:0] MUX8_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX8_io_outputs_0; // @[TopModule.scala 199:48]
  wire [3:0] MUX9_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX9_io_outputs_0; // @[TopModule.scala 199:48]
  wire [3:0] MUX10_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX10_io_outputs_0; // @[TopModule.scala 199:48]
  wire [3:0] MUX11_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX11_io_outputs_0; // @[TopModule.scala 199:48]
  wire [3:0] MUX12_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX12_io_outputs_0; // @[TopModule.scala 199:48]
  wire [3:0] MUX13_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX13_io_outputs_0; // @[TopModule.scala 199:48]
  wire [3:0] MUX14_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX14_io_outputs_0; // @[TopModule.scala 199:48]
  wire [3:0] MUX15_io_cfg; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_0; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_1; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_2; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_3; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_4; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_5; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_6; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_7; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_inputs_8; // @[TopModule.scala 199:48]
  wire [32:0] MUX15_io_outputs_0; // @[TopModule.scala 199:48]
  wire  CfgMem_clock; // @[TopModule.scala 232:29]
  wire  CfgMem_reset; // @[TopModule.scala 232:29]
  wire  CfgMem_io_cfgEn; // @[TopModule.scala 232:29]
  wire  CfgMem_io_cfgAddr; // @[TopModule.scala 232:29]
  wire [31:0] CfgMem_io_cfgData; // @[TopModule.scala 232:29]
  wire [63:0] CfgMem_io_cfgOut; // @[TopModule.scala 232:29]
  MUX0_2 MUX0 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX0_io_cfg),
    .io_inputs_0(MUX0_io_inputs_0),
    .io_inputs_1(MUX0_io_inputs_1),
    .io_inputs_2(MUX0_io_inputs_2),
    .io_inputs_3(MUX0_io_inputs_3),
    .io_inputs_4(MUX0_io_inputs_4),
    .io_inputs_5(MUX0_io_inputs_5),
    .io_inputs_6(MUX0_io_inputs_6),
    .io_inputs_7(MUX0_io_inputs_7),
    .io_inputs_8(MUX0_io_inputs_8),
    .io_outputs_0(MUX0_io_outputs_0)
  );
  MUX0_2 MUX1 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX1_io_cfg),
    .io_inputs_0(MUX1_io_inputs_0),
    .io_inputs_1(MUX1_io_inputs_1),
    .io_inputs_2(MUX1_io_inputs_2),
    .io_inputs_3(MUX1_io_inputs_3),
    .io_inputs_4(MUX1_io_inputs_4),
    .io_inputs_5(MUX1_io_inputs_5),
    .io_inputs_6(MUX1_io_inputs_6),
    .io_inputs_7(MUX1_io_inputs_7),
    .io_inputs_8(MUX1_io_inputs_8),
    .io_outputs_0(MUX1_io_outputs_0)
  );
  MUX0_2 MUX2 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX2_io_cfg),
    .io_inputs_0(MUX2_io_inputs_0),
    .io_inputs_1(MUX2_io_inputs_1),
    .io_inputs_2(MUX2_io_inputs_2),
    .io_inputs_3(MUX2_io_inputs_3),
    .io_inputs_4(MUX2_io_inputs_4),
    .io_inputs_5(MUX2_io_inputs_5),
    .io_inputs_6(MUX2_io_inputs_6),
    .io_inputs_7(MUX2_io_inputs_7),
    .io_inputs_8(MUX2_io_inputs_8),
    .io_outputs_0(MUX2_io_outputs_0)
  );
  MUX0_2 MUX3 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX3_io_cfg),
    .io_inputs_0(MUX3_io_inputs_0),
    .io_inputs_1(MUX3_io_inputs_1),
    .io_inputs_2(MUX3_io_inputs_2),
    .io_inputs_3(MUX3_io_inputs_3),
    .io_inputs_4(MUX3_io_inputs_4),
    .io_inputs_5(MUX3_io_inputs_5),
    .io_inputs_6(MUX3_io_inputs_6),
    .io_inputs_7(MUX3_io_inputs_7),
    .io_inputs_8(MUX3_io_inputs_8),
    .io_outputs_0(MUX3_io_outputs_0)
  );
  MUX0_2 MUX4 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX4_io_cfg),
    .io_inputs_0(MUX4_io_inputs_0),
    .io_inputs_1(MUX4_io_inputs_1),
    .io_inputs_2(MUX4_io_inputs_2),
    .io_inputs_3(MUX4_io_inputs_3),
    .io_inputs_4(MUX4_io_inputs_4),
    .io_inputs_5(MUX4_io_inputs_5),
    .io_inputs_6(MUX4_io_inputs_6),
    .io_inputs_7(MUX4_io_inputs_7),
    .io_inputs_8(MUX4_io_inputs_8),
    .io_outputs_0(MUX4_io_outputs_0)
  );
  MUX0_2 MUX5 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX5_io_cfg),
    .io_inputs_0(MUX5_io_inputs_0),
    .io_inputs_1(MUX5_io_inputs_1),
    .io_inputs_2(MUX5_io_inputs_2),
    .io_inputs_3(MUX5_io_inputs_3),
    .io_inputs_4(MUX5_io_inputs_4),
    .io_inputs_5(MUX5_io_inputs_5),
    .io_inputs_6(MUX5_io_inputs_6),
    .io_inputs_7(MUX5_io_inputs_7),
    .io_inputs_8(MUX5_io_inputs_8),
    .io_outputs_0(MUX5_io_outputs_0)
  );
  MUX0_2 MUX6 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX6_io_cfg),
    .io_inputs_0(MUX6_io_inputs_0),
    .io_inputs_1(MUX6_io_inputs_1),
    .io_inputs_2(MUX6_io_inputs_2),
    .io_inputs_3(MUX6_io_inputs_3),
    .io_inputs_4(MUX6_io_inputs_4),
    .io_inputs_5(MUX6_io_inputs_5),
    .io_inputs_6(MUX6_io_inputs_6),
    .io_inputs_7(MUX6_io_inputs_7),
    .io_inputs_8(MUX6_io_inputs_8),
    .io_outputs_0(MUX6_io_outputs_0)
  );
  MUX0_2 MUX7 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX7_io_cfg),
    .io_inputs_0(MUX7_io_inputs_0),
    .io_inputs_1(MUX7_io_inputs_1),
    .io_inputs_2(MUX7_io_inputs_2),
    .io_inputs_3(MUX7_io_inputs_3),
    .io_inputs_4(MUX7_io_inputs_4),
    .io_inputs_5(MUX7_io_inputs_5),
    .io_inputs_6(MUX7_io_inputs_6),
    .io_inputs_7(MUX7_io_inputs_7),
    .io_inputs_8(MUX7_io_inputs_8),
    .io_outputs_0(MUX7_io_outputs_0)
  );
  MUX0_2 MUX8 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX8_io_cfg),
    .io_inputs_0(MUX8_io_inputs_0),
    .io_inputs_1(MUX8_io_inputs_1),
    .io_inputs_2(MUX8_io_inputs_2),
    .io_inputs_3(MUX8_io_inputs_3),
    .io_inputs_4(MUX8_io_inputs_4),
    .io_inputs_5(MUX8_io_inputs_5),
    .io_inputs_6(MUX8_io_inputs_6),
    .io_inputs_7(MUX8_io_inputs_7),
    .io_inputs_8(MUX8_io_inputs_8),
    .io_outputs_0(MUX8_io_outputs_0)
  );
  MUX0_2 MUX9 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX9_io_cfg),
    .io_inputs_0(MUX9_io_inputs_0),
    .io_inputs_1(MUX9_io_inputs_1),
    .io_inputs_2(MUX9_io_inputs_2),
    .io_inputs_3(MUX9_io_inputs_3),
    .io_inputs_4(MUX9_io_inputs_4),
    .io_inputs_5(MUX9_io_inputs_5),
    .io_inputs_6(MUX9_io_inputs_6),
    .io_inputs_7(MUX9_io_inputs_7),
    .io_inputs_8(MUX9_io_inputs_8),
    .io_outputs_0(MUX9_io_outputs_0)
  );
  MUX0_2 MUX10 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX10_io_cfg),
    .io_inputs_0(MUX10_io_inputs_0),
    .io_inputs_1(MUX10_io_inputs_1),
    .io_inputs_2(MUX10_io_inputs_2),
    .io_inputs_3(MUX10_io_inputs_3),
    .io_inputs_4(MUX10_io_inputs_4),
    .io_inputs_5(MUX10_io_inputs_5),
    .io_inputs_6(MUX10_io_inputs_6),
    .io_inputs_7(MUX10_io_inputs_7),
    .io_inputs_8(MUX10_io_inputs_8),
    .io_outputs_0(MUX10_io_outputs_0)
  );
  MUX0_2 MUX11 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX11_io_cfg),
    .io_inputs_0(MUX11_io_inputs_0),
    .io_inputs_1(MUX11_io_inputs_1),
    .io_inputs_2(MUX11_io_inputs_2),
    .io_inputs_3(MUX11_io_inputs_3),
    .io_inputs_4(MUX11_io_inputs_4),
    .io_inputs_5(MUX11_io_inputs_5),
    .io_inputs_6(MUX11_io_inputs_6),
    .io_inputs_7(MUX11_io_inputs_7),
    .io_inputs_8(MUX11_io_inputs_8),
    .io_outputs_0(MUX11_io_outputs_0)
  );
  MUX0_2 MUX12 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX12_io_cfg),
    .io_inputs_0(MUX12_io_inputs_0),
    .io_inputs_1(MUX12_io_inputs_1),
    .io_inputs_2(MUX12_io_inputs_2),
    .io_inputs_3(MUX12_io_inputs_3),
    .io_inputs_4(MUX12_io_inputs_4),
    .io_inputs_5(MUX12_io_inputs_5),
    .io_inputs_6(MUX12_io_inputs_6),
    .io_inputs_7(MUX12_io_inputs_7),
    .io_inputs_8(MUX12_io_inputs_8),
    .io_outputs_0(MUX12_io_outputs_0)
  );
  MUX0_2 MUX13 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX13_io_cfg),
    .io_inputs_0(MUX13_io_inputs_0),
    .io_inputs_1(MUX13_io_inputs_1),
    .io_inputs_2(MUX13_io_inputs_2),
    .io_inputs_3(MUX13_io_inputs_3),
    .io_inputs_4(MUX13_io_inputs_4),
    .io_inputs_5(MUX13_io_inputs_5),
    .io_inputs_6(MUX13_io_inputs_6),
    .io_inputs_7(MUX13_io_inputs_7),
    .io_inputs_8(MUX13_io_inputs_8),
    .io_outputs_0(MUX13_io_outputs_0)
  );
  MUX0_2 MUX14 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX14_io_cfg),
    .io_inputs_0(MUX14_io_inputs_0),
    .io_inputs_1(MUX14_io_inputs_1),
    .io_inputs_2(MUX14_io_inputs_2),
    .io_inputs_3(MUX14_io_inputs_3),
    .io_inputs_4(MUX14_io_inputs_4),
    .io_inputs_5(MUX14_io_inputs_5),
    .io_inputs_6(MUX14_io_inputs_6),
    .io_inputs_7(MUX14_io_inputs_7),
    .io_inputs_8(MUX14_io_inputs_8),
    .io_outputs_0(MUX14_io_outputs_0)
  );
  MUX0_2 MUX15 ( // @[TopModule.scala 199:48]
    .io_cfg(MUX15_io_cfg),
    .io_inputs_0(MUX15_io_inputs_0),
    .io_inputs_1(MUX15_io_inputs_1),
    .io_inputs_2(MUX15_io_inputs_2),
    .io_inputs_3(MUX15_io_inputs_3),
    .io_inputs_4(MUX15_io_inputs_4),
    .io_inputs_5(MUX15_io_inputs_5),
    .io_inputs_6(MUX15_io_inputs_6),
    .io_inputs_7(MUX15_io_inputs_7),
    .io_inputs_8(MUX15_io_inputs_8),
    .io_outputs_0(MUX15_io_outputs_0)
  );
  CfgMem_18 CfgMem ( // @[TopModule.scala 232:29]
    .clock(CfgMem_clock),
    .reset(CfgMem_reset),
    .io_cfgEn(CfgMem_io_cfgEn),
    .io_cfgAddr(CfgMem_io_cfgAddr),
    .io_cfgData(CfgMem_io_cfgData),
    .io_cfgOut(CfgMem_io_cfgOut)
  );
  assign io_outputs_0 = MUX0_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_1 = MUX1_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_2 = MUX2_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_3 = MUX3_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_4 = MUX4_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_5 = MUX5_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_6 = MUX6_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_7 = MUX7_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_8 = MUX8_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_9 = MUX9_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_10 = MUX10_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_11 = MUX11_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_12 = MUX12_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_13 = MUX13_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_14 = MUX14_io_outputs_0; // @[TopModule.scala 392:22]
  assign io_outputs_15 = MUX15_io_outputs_0; // @[TopModule.scala 392:22]
  assign MUX0_io_cfg = CfgMem_io_cfgOut[3:0]; // @[TopModule.scala 261:98]
  assign MUX0_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX0_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX1_io_cfg = CfgMem_io_cfgOut[7:4]; // @[TopModule.scala 261:98]
  assign MUX1_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX1_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX2_io_cfg = CfgMem_io_cfgOut[11:8]; // @[TopModule.scala 261:98]
  assign MUX2_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX2_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX3_io_cfg = CfgMem_io_cfgOut[15:12]; // @[TopModule.scala 261:98]
  assign MUX3_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX3_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX4_io_cfg = CfgMem_io_cfgOut[19:16]; // @[TopModule.scala 261:98]
  assign MUX4_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX4_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX5_io_cfg = CfgMem_io_cfgOut[23:20]; // @[TopModule.scala 261:98]
  assign MUX5_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX5_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX6_io_cfg = CfgMem_io_cfgOut[27:24]; // @[TopModule.scala 261:98]
  assign MUX6_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX6_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX7_io_cfg = CfgMem_io_cfgOut[31:28]; // @[TopModule.scala 261:98]
  assign MUX7_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX7_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX8_io_cfg = CfgMem_io_cfgOut[35:32]; // @[TopModule.scala 261:98]
  assign MUX8_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX8_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX9_io_cfg = CfgMem_io_cfgOut[39:36]; // @[TopModule.scala 261:98]
  assign MUX9_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX9_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX10_io_cfg = CfgMem_io_cfgOut[43:40]; // @[TopModule.scala 261:98]
  assign MUX10_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX10_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX11_io_cfg = CfgMem_io_cfgOut[47:44]; // @[TopModule.scala 261:98]
  assign MUX11_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX11_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX12_io_cfg = CfgMem_io_cfgOut[51:48]; // @[TopModule.scala 261:98]
  assign MUX12_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX12_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX13_io_cfg = CfgMem_io_cfgOut[55:52]; // @[TopModule.scala 261:98]
  assign MUX13_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX13_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX14_io_cfg = CfgMem_io_cfgOut[59:56]; // @[TopModule.scala 261:98]
  assign MUX14_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX14_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign MUX15_io_cfg = CfgMem_io_cfgOut[63:60]; // @[TopModule.scala 261:98]
  assign MUX15_io_inputs_0 = io_inputs_0; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_1 = io_inputs_1; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_2 = io_inputs_2; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_3 = io_inputs_3; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_4 = io_inputs_4; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_5 = io_inputs_5; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_6 = io_inputs_6; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_7 = io_inputs_7; // @[TopModule.scala 392:22]
  assign MUX15_io_inputs_8 = io_inputs_8; // @[TopModule.scala 392:22]
  assign CfgMem_clock = clock;
  assign CfgMem_reset = reset;
  assign CfgMem_io_cfgEn = io_cfgEn; // @[TopModule.scala 239:34]
  assign CfgMem_io_cfgAddr = io_cfgAddr[0]; // @[TopModule.scala 244:30]
  assign CfgMem_io_cfgData = io_cfgData; // @[TopModule.scala 248:28]
endmodule
module IB0(
  input  [32:0] io_inputs_0,
  output [32:0] io_outputs_0
);
  assign io_outputs_0 = io_inputs_0; // @[IOB.scala 15:17]
endmodule
module OB0(
  input         io_cfg,
  input  [32:0] io_inputs_0,
  output [32:0] io_outputs_0
);
  wire  _T = ~io_cfg; // @[Mux.scala 80:60]
  assign io_outputs_0 = _T ? io_inputs_0 : 33'h0; // @[IOB.scala 31:19]
endmodule
module CfgMem_19(
  input         clock,
  input         reset,
  input         io_cfgEn,
  input  [31:0] io_cfgData,
  output [15:0] io_cfgOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] outWire_0; // @[Reg.scala 27:20]
  assign io_cfgOut = outWire_0[15:0]; // @[CfgMem.scala 22:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  outWire_0 = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      outWire_0 <= 32'h0;
    end else if (io_cfgEn) begin
      outWire_0 <= io_cfgData;
    end
  end
endmodule
module CGRAJ(
  input         clock,
  input         reset,
  input         io_cfgEn,
  input  [8:0]  io_cfgAddr,
  input  [31:0] io_cfgData,
  input  [32:0] io_inputs_0,
  input  [32:0] io_inputs_1,
  input  [32:0] io_inputs_2,
  input  [32:0] io_inputs_3,
  input  [32:0] io_inputs_4,
  input  [32:0] io_inputs_5,
  input  [32:0] io_inputs_6,
  input  [32:0] io_inputs_7,
  input  [32:0] io_inputs_8,
  input  [32:0] io_inputs_9,
  input  [32:0] io_inputs_10,
  input  [32:0] io_inputs_11,
  input  [32:0] io_inputs_12,
  input  [32:0] io_inputs_13,
  input  [32:0] io_inputs_14,
  input  [32:0] io_inputs_15,
  output [32:0] io_outputs_0,
  output [32:0] io_outputs_1,
  output [32:0] io_outputs_2,
  output [32:0] io_outputs_3,
  output [32:0] io_outputs_4,
  output [32:0] io_outputs_5,
  output [32:0] io_outputs_6,
  output [32:0] io_outputs_7,
  output [32:0] io_outputs_8,
  output [32:0] io_outputs_9,
  output [32:0] io_outputs_10,
  output [32:0] io_outputs_11,
  output [32:0] io_outputs_12,
  output [32:0] io_outputs_13,
  output [32:0] io_outputs_14,
  output [32:0] io_outputs_15
);
  wire  PE0_clock; // @[TopModule.scala 157:31]
  wire  PE0_reset; // @[TopModule.scala 157:31]
  wire  PE0_io_cfgEn; // @[TopModule.scala 157:31]
  wire [31:0] PE0_io_cfgData; // @[TopModule.scala 157:31]
  wire [32:0] PE0_io_inputs_0; // @[TopModule.scala 157:31]
  wire [32:0] PE0_io_inputs_1; // @[TopModule.scala 157:31]
  wire [32:0] PE0_io_outputs_0; // @[TopModule.scala 157:31]
  wire  PE1_clock; // @[TopModule.scala 157:31]
  wire  PE1_reset; // @[TopModule.scala 157:31]
  wire  PE1_io_cfgEn; // @[TopModule.scala 157:31]
  wire [31:0] PE1_io_cfgData; // @[TopModule.scala 157:31]
  wire [32:0] PE1_io_inputs_0; // @[TopModule.scala 157:31]
  wire [32:0] PE1_io_inputs_1; // @[TopModule.scala 157:31]
  wire [32:0] PE1_io_outputs_0; // @[TopModule.scala 157:31]
  wire  PE2_clock; // @[TopModule.scala 157:31]
  wire  PE2_reset; // @[TopModule.scala 157:31]
  wire  PE2_io_cfgEn; // @[TopModule.scala 157:31]
  wire [31:0] PE2_io_cfgData; // @[TopModule.scala 157:31]
  wire [32:0] PE2_io_inputs_0; // @[TopModule.scala 157:31]
  wire [32:0] PE2_io_inputs_1; // @[TopModule.scala 157:31]
  wire [32:0] PE2_io_outputs_0; // @[TopModule.scala 157:31]
  wire  PE3_clock; // @[TopModule.scala 157:31]
  wire  PE3_reset; // @[TopModule.scala 157:31]
  wire  PE3_io_cfgEn; // @[TopModule.scala 157:31]
  wire [31:0] PE3_io_cfgData; // @[TopModule.scala 157:31]
  wire [32:0] PE3_io_inputs_0; // @[TopModule.scala 157:31]
  wire [32:0] PE3_io_inputs_1; // @[TopModule.scala 157:31]
  wire [32:0] PE3_io_outputs_0; // @[TopModule.scala 157:31]
  wire  PE4_clock; // @[TopModule.scala 157:31]
  wire  PE4_reset; // @[TopModule.scala 157:31]
  wire  PE4_io_cfgEn; // @[TopModule.scala 157:31]
  wire [31:0] PE4_io_cfgData; // @[TopModule.scala 157:31]
  wire [32:0] PE4_io_inputs_0; // @[TopModule.scala 157:31]
  wire [32:0] PE4_io_inputs_1; // @[TopModule.scala 157:31]
  wire [32:0] PE4_io_outputs_0; // @[TopModule.scala 157:31]
  wire  PE5_clock; // @[TopModule.scala 157:31]
  wire  PE5_reset; // @[TopModule.scala 157:31]
  wire  PE5_io_cfgEn; // @[TopModule.scala 157:31]
  wire [31:0] PE5_io_cfgData; // @[TopModule.scala 157:31]
  wire [32:0] PE5_io_inputs_0; // @[TopModule.scala 157:31]
  wire [32:0] PE5_io_inputs_1; // @[TopModule.scala 157:31]
  wire [32:0] PE5_io_outputs_0; // @[TopModule.scala 157:31]
  wire  PE6_clock; // @[TopModule.scala 157:31]
  wire  PE6_reset; // @[TopModule.scala 157:31]
  wire  PE6_io_cfgEn; // @[TopModule.scala 157:31]
  wire [31:0] PE6_io_cfgData; // @[TopModule.scala 157:31]
  wire [32:0] PE6_io_inputs_0; // @[TopModule.scala 157:31]
  wire [32:0] PE6_io_inputs_1; // @[TopModule.scala 157:31]
  wire [32:0] PE6_io_outputs_0; // @[TopModule.scala 157:31]
  wire  PE7_clock; // @[TopModule.scala 157:31]
  wire  PE7_reset; // @[TopModule.scala 157:31]
  wire  PE7_io_cfgEn; // @[TopModule.scala 157:31]
  wire [31:0] PE7_io_cfgData; // @[TopModule.scala 157:31]
  wire [32:0] PE7_io_inputs_0; // @[TopModule.scala 157:31]
  wire [32:0] PE7_io_inputs_1; // @[TopModule.scala 157:31]
  wire [32:0] PE7_io_outputs_0; // @[TopModule.scala 157:31]
  wire  PE8_clock; // @[TopModule.scala 157:31]
  wire  PE8_reset; // @[TopModule.scala 157:31]
  wire  PE8_io_cfgEn; // @[TopModule.scala 157:31]
  wire [31:0] PE8_io_cfgData; // @[TopModule.scala 157:31]
  wire [32:0] PE8_io_inputs_0; // @[TopModule.scala 157:31]
  wire [32:0] PE8_io_inputs_1; // @[TopModule.scala 157:31]
  wire [32:0] PE8_io_outputs_0; // @[TopModule.scala 157:31]
  wire [32:0] dpicDebug_in; // @[TopModule.scala 165:33]
  wire  PE9_clock; // @[TopModule.scala 157:31]
  wire  PE9_reset; // @[TopModule.scala 157:31]
  wire  PE9_io_cfgEn; // @[TopModule.scala 157:31]
  wire [31:0] PE9_io_cfgData; // @[TopModule.scala 157:31]
  wire [32:0] PE9_io_inputs_0; // @[TopModule.scala 157:31]
  wire [32:0] PE9_io_inputs_1; // @[TopModule.scala 157:31]
  wire [32:0] PE9_io_outputs_0; // @[TopModule.scala 157:31]
  wire  PE10_clock; // @[TopModule.scala 157:31]
  wire  PE10_reset; // @[TopModule.scala 157:31]
  wire  PE10_io_cfgEn; // @[TopModule.scala 157:31]
  wire [31:0] PE10_io_cfgData; // @[TopModule.scala 157:31]
  wire [32:0] PE10_io_inputs_0; // @[TopModule.scala 157:31]
  wire [32:0] PE10_io_inputs_1; // @[TopModule.scala 157:31]
  wire [32:0] PE10_io_outputs_0; // @[TopModule.scala 157:31]
  wire  PE11_clock; // @[TopModule.scala 157:31]
  wire  PE11_reset; // @[TopModule.scala 157:31]
  wire  PE11_io_cfgEn; // @[TopModule.scala 157:31]
  wire [31:0] PE11_io_cfgData; // @[TopModule.scala 157:31]
  wire [32:0] PE11_io_inputs_0; // @[TopModule.scala 157:31]
  wire [32:0] PE11_io_inputs_1; // @[TopModule.scala 157:31]
  wire [32:0] PE11_io_outputs_0; // @[TopModule.scala 157:31]
  wire  PE12_clock; // @[TopModule.scala 157:31]
  wire  PE12_reset; // @[TopModule.scala 157:31]
  wire  PE12_io_cfgEn; // @[TopModule.scala 157:31]
  wire [31:0] PE12_io_cfgData; // @[TopModule.scala 157:31]
  wire [32:0] PE12_io_inputs_0; // @[TopModule.scala 157:31]
  wire [32:0] PE12_io_inputs_1; // @[TopModule.scala 157:31]
  wire [32:0] PE12_io_outputs_0; // @[TopModule.scala 157:31]
  wire  PE13_clock; // @[TopModule.scala 157:31]
  wire  PE13_reset; // @[TopModule.scala 157:31]
  wire  PE13_io_cfgEn; // @[TopModule.scala 157:31]
  wire [31:0] PE13_io_cfgData; // @[TopModule.scala 157:31]
  wire [32:0] PE13_io_inputs_0; // @[TopModule.scala 157:31]
  wire [32:0] PE13_io_inputs_1; // @[TopModule.scala 157:31]
  wire [32:0] PE13_io_outputs_0; // @[TopModule.scala 157:31]
  wire  PE14_clock; // @[TopModule.scala 157:31]
  wire  PE14_reset; // @[TopModule.scala 157:31]
  wire  PE14_io_cfgEn; // @[TopModule.scala 157:31]
  wire [31:0] PE14_io_cfgData; // @[TopModule.scala 157:31]
  wire [32:0] PE14_io_inputs_0; // @[TopModule.scala 157:31]
  wire [32:0] PE14_io_inputs_1; // @[TopModule.scala 157:31]
  wire [32:0] PE14_io_outputs_0; // @[TopModule.scala 157:31]
  wire  PE15_clock; // @[TopModule.scala 157:31]
  wire  PE15_reset; // @[TopModule.scala 157:31]
  wire  PE15_io_cfgEn; // @[TopModule.scala 157:31]
  wire [31:0] PE15_io_cfgData; // @[TopModule.scala 157:31]
  wire [32:0] PE15_io_inputs_0; // @[TopModule.scala 157:31]
  wire [32:0] PE15_io_inputs_1; // @[TopModule.scala 157:31]
  wire [32:0] PE15_io_outputs_0; // @[TopModule.scala 157:31]
  wire  MatrixFC0_clock; // @[TopModule.scala 157:31]
  wire  MatrixFC0_reset; // @[TopModule.scala 157:31]
  wire  MatrixFC0_io_cfgEn; // @[TopModule.scala 157:31]
  wire [3:0] MatrixFC0_io_cfgAddr; // @[TopModule.scala 157:31]
  wire [31:0] MatrixFC0_io_cfgData; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_inputs_0; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_inputs_1; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_inputs_2; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_inputs_3; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_inputs_4; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_inputs_5; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_inputs_6; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_inputs_7; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_inputs_8; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_inputs_9; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_inputs_10; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_inputs_11; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_inputs_12; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_inputs_13; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_inputs_14; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_inputs_15; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_inputs_16; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_outputs_0; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_outputs_1; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_outputs_2; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_outputs_3; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_outputs_4; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_outputs_5; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_outputs_6; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_outputs_7; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_outputs_8; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_outputs_9; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_outputs_10; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_outputs_11; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_outputs_12; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_outputs_13; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_outputs_14; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_outputs_15; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC0_io_outputs_16; // @[TopModule.scala 157:31]
  wire  MatrixFC1_clock; // @[TopModule.scala 157:31]
  wire  MatrixFC1_reset; // @[TopModule.scala 157:31]
  wire  MatrixFC1_io_cfgEn; // @[TopModule.scala 157:31]
  wire [3:0] MatrixFC1_io_cfgAddr; // @[TopModule.scala 157:31]
  wire [31:0] MatrixFC1_io_cfgData; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_0; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_1; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_2; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_3; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_4; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_5; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_6; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_7; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_8; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_9; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_10; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_11; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_12; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_13; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_14; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_15; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_16; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_17; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_18; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_19; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_20; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_21; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_22; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_inputs_23; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_outputs_0; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_outputs_1; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_outputs_2; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_outputs_3; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_outputs_4; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_outputs_5; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_outputs_6; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_outputs_7; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_outputs_8; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_outputs_9; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_outputs_10; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_outputs_11; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_outputs_12; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_outputs_13; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_outputs_14; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_outputs_15; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC1_io_outputs_16; // @[TopModule.scala 157:31]
  wire  MatrixFC2_clock; // @[TopModule.scala 157:31]
  wire  MatrixFC2_reset; // @[TopModule.scala 157:31]
  wire  MatrixFC2_io_cfgEn; // @[TopModule.scala 157:31]
  wire [3:0] MatrixFC2_io_cfgAddr; // @[TopModule.scala 157:31]
  wire [31:0] MatrixFC2_io_cfgData; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_inputs_0; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_inputs_1; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_inputs_2; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_inputs_3; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_inputs_4; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_inputs_5; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_inputs_6; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_inputs_7; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_inputs_8; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_outputs_0; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_outputs_1; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_outputs_2; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_outputs_3; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_outputs_4; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_outputs_5; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_outputs_6; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_outputs_7; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_outputs_8; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_outputs_9; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_outputs_10; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_outputs_11; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_outputs_12; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_outputs_13; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_outputs_14; // @[TopModule.scala 157:31]
  wire [32:0] MatrixFC2_io_outputs_15; // @[TopModule.scala 157:31]
  wire [32:0] IB0_io_inputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB0_io_outputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB1_io_inputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB1_io_outputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB2_io_inputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB2_io_outputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB3_io_inputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB3_io_outputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB4_io_inputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB4_io_outputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB5_io_inputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB5_io_outputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB6_io_inputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB6_io_outputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB7_io_inputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB7_io_outputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB8_io_inputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB8_io_outputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB9_io_inputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB9_io_outputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB10_io_inputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB10_io_outputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB11_io_inputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB11_io_outputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB12_io_inputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB12_io_outputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB13_io_inputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB13_io_outputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB14_io_inputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB14_io_outputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB15_io_inputs_0; // @[TopModule.scala 216:48]
  wire [32:0] IB15_io_outputs_0; // @[TopModule.scala 216:48]
  wire  OB0_io_cfg; // @[TopModule.scala 220:48]
  wire [32:0] OB0_io_inputs_0; // @[TopModule.scala 220:48]
  wire [32:0] OB0_io_outputs_0; // @[TopModule.scala 220:48]
  wire  OB1_io_cfg; // @[TopModule.scala 220:48]
  wire [32:0] OB1_io_inputs_0; // @[TopModule.scala 220:48]
  wire [32:0] OB1_io_outputs_0; // @[TopModule.scala 220:48]
  wire  OB2_io_cfg; // @[TopModule.scala 220:48]
  wire [32:0] OB2_io_inputs_0; // @[TopModule.scala 220:48]
  wire [32:0] OB2_io_outputs_0; // @[TopModule.scala 220:48]
  wire  OB3_io_cfg; // @[TopModule.scala 220:48]
  wire [32:0] OB3_io_inputs_0; // @[TopModule.scala 220:48]
  wire [32:0] OB3_io_outputs_0; // @[TopModule.scala 220:48]
  wire  OB4_io_cfg; // @[TopModule.scala 220:48]
  wire [32:0] OB4_io_inputs_0; // @[TopModule.scala 220:48]
  wire [32:0] OB4_io_outputs_0; // @[TopModule.scala 220:48]
  wire  OB5_io_cfg; // @[TopModule.scala 220:48]
  wire [32:0] OB5_io_inputs_0; // @[TopModule.scala 220:48]
  wire [32:0] OB5_io_outputs_0; // @[TopModule.scala 220:48]
  wire  OB6_io_cfg; // @[TopModule.scala 220:48]
  wire [32:0] OB6_io_inputs_0; // @[TopModule.scala 220:48]
  wire [32:0] OB6_io_outputs_0; // @[TopModule.scala 220:48]
  wire  OB7_io_cfg; // @[TopModule.scala 220:48]
  wire [32:0] OB7_io_inputs_0; // @[TopModule.scala 220:48]
  wire [32:0] OB7_io_outputs_0; // @[TopModule.scala 220:48]
  wire  OB8_io_cfg; // @[TopModule.scala 220:48]
  wire [32:0] OB8_io_inputs_0; // @[TopModule.scala 220:48]
  wire [32:0] OB8_io_outputs_0; // @[TopModule.scala 220:48]
  wire  OB9_io_cfg; // @[TopModule.scala 220:48]
  wire [32:0] OB9_io_inputs_0; // @[TopModule.scala 220:48]
  wire [32:0] OB9_io_outputs_0; // @[TopModule.scala 220:48]
  wire  OB10_io_cfg; // @[TopModule.scala 220:48]
  wire [32:0] OB10_io_inputs_0; // @[TopModule.scala 220:48]
  wire [32:0] OB10_io_outputs_0; // @[TopModule.scala 220:48]
  wire  OB11_io_cfg; // @[TopModule.scala 220:48]
  wire [32:0] OB11_io_inputs_0; // @[TopModule.scala 220:48]
  wire [32:0] OB11_io_outputs_0; // @[TopModule.scala 220:48]
  wire  OB12_io_cfg; // @[TopModule.scala 220:48]
  wire [32:0] OB12_io_inputs_0; // @[TopModule.scala 220:48]
  wire [32:0] OB12_io_outputs_0; // @[TopModule.scala 220:48]
  wire  OB13_io_cfg; // @[TopModule.scala 220:48]
  wire [32:0] OB13_io_inputs_0; // @[TopModule.scala 220:48]
  wire [32:0] OB13_io_outputs_0; // @[TopModule.scala 220:48]
  wire  OB14_io_cfg; // @[TopModule.scala 220:48]
  wire [32:0] OB14_io_inputs_0; // @[TopModule.scala 220:48]
  wire [32:0] OB14_io_outputs_0; // @[TopModule.scala 220:48]
  wire  OB15_io_cfg; // @[TopModule.scala 220:48]
  wire [32:0] OB15_io_inputs_0; // @[TopModule.scala 220:48]
  wire [32:0] OB15_io_outputs_0; // @[TopModule.scala 220:48]
  wire  CfgMem_clock; // @[TopModule.scala 232:29]
  wire  CfgMem_reset; // @[TopModule.scala 232:29]
  wire  CfgMem_io_cfgEn; // @[TopModule.scala 232:29]
  wire [31:0] CfgMem_io_cfgData; // @[TopModule.scala 232:29]
  wire [15:0] CfgMem_io_cfgOut; // @[TopModule.scala 232:29]
  wire [32:0] dpicCGRA_ins_0; // @[TopModule.scala 292:27]
  wire [32:0] dpicCGRA_ins_1; // @[TopModule.scala 292:27]
  wire [32:0] dpicCGRA_ins_2; // @[TopModule.scala 292:27]
  wire [32:0] dpicCGRA_ins_3; // @[TopModule.scala 292:27]
  wire [32:0] dpicCGRA_ins_4; // @[TopModule.scala 292:27]
  wire [32:0] dpicCGRA_ins_5; // @[TopModule.scala 292:27]
  wire [32:0] dpicCGRA_ins_6; // @[TopModule.scala 292:27]
  wire [32:0] dpicCGRA_ins_7; // @[TopModule.scala 292:27]
  wire [32:0] dpicCGRA_ins_8; // @[TopModule.scala 292:27]
  wire [32:0] dpicCGRA_ins_9; // @[TopModule.scala 292:27]
  wire [32:0] dpicCGRA_ins_10; // @[TopModule.scala 292:27]
  wire [32:0] dpicCGRA_ins_11; // @[TopModule.scala 292:27]
  wire [32:0] dpicCGRA_ins_12; // @[TopModule.scala 292:27]
  wire [32:0] dpicCGRA_ins_13; // @[TopModule.scala 292:27]
  wire [32:0] dpicCGRA_ins_14; // @[TopModule.scala 292:27]
  wire [32:0] dpicCGRA_ins_15; // @[TopModule.scala 292:27]
  wire  _T_1 = io_cfgAddr[8:4] == 5'h1; // @[TopModule.scala 159:106]
  wire  _T_4 = io_cfgAddr[8:4] == 5'h2; // @[TopModule.scala 159:106]
  wire  _T_7 = io_cfgAddr[8:4] == 5'h3; // @[TopModule.scala 159:106]
  wire  _T_10 = io_cfgAddr[8:4] == 5'h4; // @[TopModule.scala 159:106]
  wire  _T_13 = io_cfgAddr[8:4] == 5'h5; // @[TopModule.scala 159:106]
  wire  _T_16 = io_cfgAddr[8:4] == 5'h6; // @[TopModule.scala 159:106]
  wire  _T_19 = io_cfgAddr[8:4] == 5'h7; // @[TopModule.scala 159:106]
  wire  _T_22 = io_cfgAddr[8:4] == 5'h8; // @[TopModule.scala 159:106]
  wire  _T_25 = io_cfgAddr[8:4] == 5'h9; // @[TopModule.scala 159:106]
  wire  _T_28 = io_cfgAddr[8:4] == 5'ha; // @[TopModule.scala 159:106]
  wire  _T_31 = io_cfgAddr[8:4] == 5'hb; // @[TopModule.scala 159:106]
  wire  _T_34 = io_cfgAddr[8:4] == 5'hc; // @[TopModule.scala 159:106]
  wire  _T_37 = io_cfgAddr[8:4] == 5'hd; // @[TopModule.scala 159:106]
  wire  _T_40 = io_cfgAddr[8:4] == 5'he; // @[TopModule.scala 159:106]
  wire  _T_43 = io_cfgAddr[8:4] == 5'hf; // @[TopModule.scala 159:106]
  wire  _T_46 = io_cfgAddr[8:4] == 5'h10; // @[TopModule.scala 159:106]
  wire  _T_49 = io_cfgAddr[8:4] == 5'h11; // @[TopModule.scala 159:106]
  wire  _T_52 = io_cfgAddr[8:4] == 5'h12; // @[TopModule.scala 159:106]
  wire  _T_55 = io_cfgAddr[8:4] == 5'h13; // @[TopModule.scala 159:106]
  wire  _T_58 = io_cfgAddr[8:4] == 5'h0; // @[TopModule.scala 241:109]
  PE0 PE0 ( // @[TopModule.scala 157:31]
    .clock(PE0_clock),
    .reset(PE0_reset),
    .io_cfgEn(PE0_io_cfgEn),
    .io_cfgData(PE0_io_cfgData),
    .io_inputs_0(PE0_io_inputs_0),
    .io_inputs_1(PE0_io_inputs_1),
    .io_outputs_0(PE0_io_outputs_0)
  );
  PE0 PE1 ( // @[TopModule.scala 157:31]
    .clock(PE1_clock),
    .reset(PE1_reset),
    .io_cfgEn(PE1_io_cfgEn),
    .io_cfgData(PE1_io_cfgData),
    .io_inputs_0(PE1_io_inputs_0),
    .io_inputs_1(PE1_io_inputs_1),
    .io_outputs_0(PE1_io_outputs_0)
  );
  PE0 PE2 ( // @[TopModule.scala 157:31]
    .clock(PE2_clock),
    .reset(PE2_reset),
    .io_cfgEn(PE2_io_cfgEn),
    .io_cfgData(PE2_io_cfgData),
    .io_inputs_0(PE2_io_inputs_0),
    .io_inputs_1(PE2_io_inputs_1),
    .io_outputs_0(PE2_io_outputs_0)
  );
  PE0 PE3 ( // @[TopModule.scala 157:31]
    .clock(PE3_clock),
    .reset(PE3_reset),
    .io_cfgEn(PE3_io_cfgEn),
    .io_cfgData(PE3_io_cfgData),
    .io_inputs_0(PE3_io_inputs_0),
    .io_inputs_1(PE3_io_inputs_1),
    .io_outputs_0(PE3_io_outputs_0)
  );
  PE0 PE4 ( // @[TopModule.scala 157:31]
    .clock(PE4_clock),
    .reset(PE4_reset),
    .io_cfgEn(PE4_io_cfgEn),
    .io_cfgData(PE4_io_cfgData),
    .io_inputs_0(PE4_io_inputs_0),
    .io_inputs_1(PE4_io_inputs_1),
    .io_outputs_0(PE4_io_outputs_0)
  );
  PE0 PE5 ( // @[TopModule.scala 157:31]
    .clock(PE5_clock),
    .reset(PE5_reset),
    .io_cfgEn(PE5_io_cfgEn),
    .io_cfgData(PE5_io_cfgData),
    .io_inputs_0(PE5_io_inputs_0),
    .io_inputs_1(PE5_io_inputs_1),
    .io_outputs_0(PE5_io_outputs_0)
  );
  PE0 PE6 ( // @[TopModule.scala 157:31]
    .clock(PE6_clock),
    .reset(PE6_reset),
    .io_cfgEn(PE6_io_cfgEn),
    .io_cfgData(PE6_io_cfgData),
    .io_inputs_0(PE6_io_inputs_0),
    .io_inputs_1(PE6_io_inputs_1),
    .io_outputs_0(PE6_io_outputs_0)
  );
  PE0 PE7 ( // @[TopModule.scala 157:31]
    .clock(PE7_clock),
    .reset(PE7_reset),
    .io_cfgEn(PE7_io_cfgEn),
    .io_cfgData(PE7_io_cfgData),
    .io_inputs_0(PE7_io_inputs_0),
    .io_inputs_1(PE7_io_inputs_1),
    .io_outputs_0(PE7_io_outputs_0)
  );
  PE0 PE8 ( // @[TopModule.scala 157:31]
    .clock(PE8_clock),
    .reset(PE8_reset),
    .io_cfgEn(PE8_io_cfgEn),
    .io_cfgData(PE8_io_cfgData),
    .io_inputs_0(PE8_io_inputs_0),
    .io_inputs_1(PE8_io_inputs_1),
    .io_outputs_0(PE8_io_outputs_0)
  );
  dpicDebug dpicDebug ( // @[TopModule.scala 165:33]
    .in(dpicDebug_in)
  );
  PE0 PE9 ( // @[TopModule.scala 157:31]
    .clock(PE9_clock),
    .reset(PE9_reset),
    .io_cfgEn(PE9_io_cfgEn),
    .io_cfgData(PE9_io_cfgData),
    .io_inputs_0(PE9_io_inputs_0),
    .io_inputs_1(PE9_io_inputs_1),
    .io_outputs_0(PE9_io_outputs_0)
  );
  PE0 PE10 ( // @[TopModule.scala 157:31]
    .clock(PE10_clock),
    .reset(PE10_reset),
    .io_cfgEn(PE10_io_cfgEn),
    .io_cfgData(PE10_io_cfgData),
    .io_inputs_0(PE10_io_inputs_0),
    .io_inputs_1(PE10_io_inputs_1),
    .io_outputs_0(PE10_io_outputs_0)
  );
  PE0 PE11 ( // @[TopModule.scala 157:31]
    .clock(PE11_clock),
    .reset(PE11_reset),
    .io_cfgEn(PE11_io_cfgEn),
    .io_cfgData(PE11_io_cfgData),
    .io_inputs_0(PE11_io_inputs_0),
    .io_inputs_1(PE11_io_inputs_1),
    .io_outputs_0(PE11_io_outputs_0)
  );
  PE0 PE12 ( // @[TopModule.scala 157:31]
    .clock(PE12_clock),
    .reset(PE12_reset),
    .io_cfgEn(PE12_io_cfgEn),
    .io_cfgData(PE12_io_cfgData),
    .io_inputs_0(PE12_io_inputs_0),
    .io_inputs_1(PE12_io_inputs_1),
    .io_outputs_0(PE12_io_outputs_0)
  );
  PE0 PE13 ( // @[TopModule.scala 157:31]
    .clock(PE13_clock),
    .reset(PE13_reset),
    .io_cfgEn(PE13_io_cfgEn),
    .io_cfgData(PE13_io_cfgData),
    .io_inputs_0(PE13_io_inputs_0),
    .io_inputs_1(PE13_io_inputs_1),
    .io_outputs_0(PE13_io_outputs_0)
  );
  PE0 PE14 ( // @[TopModule.scala 157:31]
    .clock(PE14_clock),
    .reset(PE14_reset),
    .io_cfgEn(PE14_io_cfgEn),
    .io_cfgData(PE14_io_cfgData),
    .io_inputs_0(PE14_io_inputs_0),
    .io_inputs_1(PE14_io_inputs_1),
    .io_outputs_0(PE14_io_outputs_0)
  );
  PE0 PE15 ( // @[TopModule.scala 157:31]
    .clock(PE15_clock),
    .reset(PE15_reset),
    .io_cfgEn(PE15_io_cfgEn),
    .io_cfgData(PE15_io_cfgData),
    .io_inputs_0(PE15_io_inputs_0),
    .io_inputs_1(PE15_io_inputs_1),
    .io_outputs_0(PE15_io_outputs_0)
  );
  matrixFCdevice0 MatrixFC0 ( // @[TopModule.scala 157:31]
    .clock(MatrixFC0_clock),
    .reset(MatrixFC0_reset),
    .io_cfgEn(MatrixFC0_io_cfgEn),
    .io_cfgAddr(MatrixFC0_io_cfgAddr),
    .io_cfgData(MatrixFC0_io_cfgData),
    .io_inputs_0(MatrixFC0_io_inputs_0),
    .io_inputs_1(MatrixFC0_io_inputs_1),
    .io_inputs_2(MatrixFC0_io_inputs_2),
    .io_inputs_3(MatrixFC0_io_inputs_3),
    .io_inputs_4(MatrixFC0_io_inputs_4),
    .io_inputs_5(MatrixFC0_io_inputs_5),
    .io_inputs_6(MatrixFC0_io_inputs_6),
    .io_inputs_7(MatrixFC0_io_inputs_7),
    .io_inputs_8(MatrixFC0_io_inputs_8),
    .io_inputs_9(MatrixFC0_io_inputs_9),
    .io_inputs_10(MatrixFC0_io_inputs_10),
    .io_inputs_11(MatrixFC0_io_inputs_11),
    .io_inputs_12(MatrixFC0_io_inputs_12),
    .io_inputs_13(MatrixFC0_io_inputs_13),
    .io_inputs_14(MatrixFC0_io_inputs_14),
    .io_inputs_15(MatrixFC0_io_inputs_15),
    .io_inputs_16(MatrixFC0_io_inputs_16),
    .io_outputs_0(MatrixFC0_io_outputs_0),
    .io_outputs_1(MatrixFC0_io_outputs_1),
    .io_outputs_2(MatrixFC0_io_outputs_2),
    .io_outputs_3(MatrixFC0_io_outputs_3),
    .io_outputs_4(MatrixFC0_io_outputs_4),
    .io_outputs_5(MatrixFC0_io_outputs_5),
    .io_outputs_6(MatrixFC0_io_outputs_6),
    .io_outputs_7(MatrixFC0_io_outputs_7),
    .io_outputs_8(MatrixFC0_io_outputs_8),
    .io_outputs_9(MatrixFC0_io_outputs_9),
    .io_outputs_10(MatrixFC0_io_outputs_10),
    .io_outputs_11(MatrixFC0_io_outputs_11),
    .io_outputs_12(MatrixFC0_io_outputs_12),
    .io_outputs_13(MatrixFC0_io_outputs_13),
    .io_outputs_14(MatrixFC0_io_outputs_14),
    .io_outputs_15(MatrixFC0_io_outputs_15),
    .io_outputs_16(MatrixFC0_io_outputs_16)
  );
  matrixFCdevice1 MatrixFC1 ( // @[TopModule.scala 157:31]
    .clock(MatrixFC1_clock),
    .reset(MatrixFC1_reset),
    .io_cfgEn(MatrixFC1_io_cfgEn),
    .io_cfgAddr(MatrixFC1_io_cfgAddr),
    .io_cfgData(MatrixFC1_io_cfgData),
    .io_inputs_0(MatrixFC1_io_inputs_0),
    .io_inputs_1(MatrixFC1_io_inputs_1),
    .io_inputs_2(MatrixFC1_io_inputs_2),
    .io_inputs_3(MatrixFC1_io_inputs_3),
    .io_inputs_4(MatrixFC1_io_inputs_4),
    .io_inputs_5(MatrixFC1_io_inputs_5),
    .io_inputs_6(MatrixFC1_io_inputs_6),
    .io_inputs_7(MatrixFC1_io_inputs_7),
    .io_inputs_8(MatrixFC1_io_inputs_8),
    .io_inputs_9(MatrixFC1_io_inputs_9),
    .io_inputs_10(MatrixFC1_io_inputs_10),
    .io_inputs_11(MatrixFC1_io_inputs_11),
    .io_inputs_12(MatrixFC1_io_inputs_12),
    .io_inputs_13(MatrixFC1_io_inputs_13),
    .io_inputs_14(MatrixFC1_io_inputs_14),
    .io_inputs_15(MatrixFC1_io_inputs_15),
    .io_inputs_16(MatrixFC1_io_inputs_16),
    .io_inputs_17(MatrixFC1_io_inputs_17),
    .io_inputs_18(MatrixFC1_io_inputs_18),
    .io_inputs_19(MatrixFC1_io_inputs_19),
    .io_inputs_20(MatrixFC1_io_inputs_20),
    .io_inputs_21(MatrixFC1_io_inputs_21),
    .io_inputs_22(MatrixFC1_io_inputs_22),
    .io_inputs_23(MatrixFC1_io_inputs_23),
    .io_outputs_0(MatrixFC1_io_outputs_0),
    .io_outputs_1(MatrixFC1_io_outputs_1),
    .io_outputs_2(MatrixFC1_io_outputs_2),
    .io_outputs_3(MatrixFC1_io_outputs_3),
    .io_outputs_4(MatrixFC1_io_outputs_4),
    .io_outputs_5(MatrixFC1_io_outputs_5),
    .io_outputs_6(MatrixFC1_io_outputs_6),
    .io_outputs_7(MatrixFC1_io_outputs_7),
    .io_outputs_8(MatrixFC1_io_outputs_8),
    .io_outputs_9(MatrixFC1_io_outputs_9),
    .io_outputs_10(MatrixFC1_io_outputs_10),
    .io_outputs_11(MatrixFC1_io_outputs_11),
    .io_outputs_12(MatrixFC1_io_outputs_12),
    .io_outputs_13(MatrixFC1_io_outputs_13),
    .io_outputs_14(MatrixFC1_io_outputs_14),
    .io_outputs_15(MatrixFC1_io_outputs_15),
    .io_outputs_16(MatrixFC1_io_outputs_16)
  );
  matrixFCdevice2 MatrixFC2 ( // @[TopModule.scala 157:31]
    .clock(MatrixFC2_clock),
    .reset(MatrixFC2_reset),
    .io_cfgEn(MatrixFC2_io_cfgEn),
    .io_cfgAddr(MatrixFC2_io_cfgAddr),
    .io_cfgData(MatrixFC2_io_cfgData),
    .io_inputs_0(MatrixFC2_io_inputs_0),
    .io_inputs_1(MatrixFC2_io_inputs_1),
    .io_inputs_2(MatrixFC2_io_inputs_2),
    .io_inputs_3(MatrixFC2_io_inputs_3),
    .io_inputs_4(MatrixFC2_io_inputs_4),
    .io_inputs_5(MatrixFC2_io_inputs_5),
    .io_inputs_6(MatrixFC2_io_inputs_6),
    .io_inputs_7(MatrixFC2_io_inputs_7),
    .io_inputs_8(MatrixFC2_io_inputs_8),
    .io_outputs_0(MatrixFC2_io_outputs_0),
    .io_outputs_1(MatrixFC2_io_outputs_1),
    .io_outputs_2(MatrixFC2_io_outputs_2),
    .io_outputs_3(MatrixFC2_io_outputs_3),
    .io_outputs_4(MatrixFC2_io_outputs_4),
    .io_outputs_5(MatrixFC2_io_outputs_5),
    .io_outputs_6(MatrixFC2_io_outputs_6),
    .io_outputs_7(MatrixFC2_io_outputs_7),
    .io_outputs_8(MatrixFC2_io_outputs_8),
    .io_outputs_9(MatrixFC2_io_outputs_9),
    .io_outputs_10(MatrixFC2_io_outputs_10),
    .io_outputs_11(MatrixFC2_io_outputs_11),
    .io_outputs_12(MatrixFC2_io_outputs_12),
    .io_outputs_13(MatrixFC2_io_outputs_13),
    .io_outputs_14(MatrixFC2_io_outputs_14),
    .io_outputs_15(MatrixFC2_io_outputs_15)
  );
  IB0 IB0 ( // @[TopModule.scala 216:48]
    .io_inputs_0(IB0_io_inputs_0),
    .io_outputs_0(IB0_io_outputs_0)
  );
  IB0 IB1 ( // @[TopModule.scala 216:48]
    .io_inputs_0(IB1_io_inputs_0),
    .io_outputs_0(IB1_io_outputs_0)
  );
  IB0 IB2 ( // @[TopModule.scala 216:48]
    .io_inputs_0(IB2_io_inputs_0),
    .io_outputs_0(IB2_io_outputs_0)
  );
  IB0 IB3 ( // @[TopModule.scala 216:48]
    .io_inputs_0(IB3_io_inputs_0),
    .io_outputs_0(IB3_io_outputs_0)
  );
  IB0 IB4 ( // @[TopModule.scala 216:48]
    .io_inputs_0(IB4_io_inputs_0),
    .io_outputs_0(IB4_io_outputs_0)
  );
  IB0 IB5 ( // @[TopModule.scala 216:48]
    .io_inputs_0(IB5_io_inputs_0),
    .io_outputs_0(IB5_io_outputs_0)
  );
  IB0 IB6 ( // @[TopModule.scala 216:48]
    .io_inputs_0(IB6_io_inputs_0),
    .io_outputs_0(IB6_io_outputs_0)
  );
  IB0 IB7 ( // @[TopModule.scala 216:48]
    .io_inputs_0(IB7_io_inputs_0),
    .io_outputs_0(IB7_io_outputs_0)
  );
  IB0 IB8 ( // @[TopModule.scala 216:48]
    .io_inputs_0(IB8_io_inputs_0),
    .io_outputs_0(IB8_io_outputs_0)
  );
  IB0 IB9 ( // @[TopModule.scala 216:48]
    .io_inputs_0(IB9_io_inputs_0),
    .io_outputs_0(IB9_io_outputs_0)
  );
  IB0 IB10 ( // @[TopModule.scala 216:48]
    .io_inputs_0(IB10_io_inputs_0),
    .io_outputs_0(IB10_io_outputs_0)
  );
  IB0 IB11 ( // @[TopModule.scala 216:48]
    .io_inputs_0(IB11_io_inputs_0),
    .io_outputs_0(IB11_io_outputs_0)
  );
  IB0 IB12 ( // @[TopModule.scala 216:48]
    .io_inputs_0(IB12_io_inputs_0),
    .io_outputs_0(IB12_io_outputs_0)
  );
  IB0 IB13 ( // @[TopModule.scala 216:48]
    .io_inputs_0(IB13_io_inputs_0),
    .io_outputs_0(IB13_io_outputs_0)
  );
  IB0 IB14 ( // @[TopModule.scala 216:48]
    .io_inputs_0(IB14_io_inputs_0),
    .io_outputs_0(IB14_io_outputs_0)
  );
  IB0 IB15 ( // @[TopModule.scala 216:48]
    .io_inputs_0(IB15_io_inputs_0),
    .io_outputs_0(IB15_io_outputs_0)
  );
  OB0 OB0 ( // @[TopModule.scala 220:48]
    .io_cfg(OB0_io_cfg),
    .io_inputs_0(OB0_io_inputs_0),
    .io_outputs_0(OB0_io_outputs_0)
  );
  OB0 OB1 ( // @[TopModule.scala 220:48]
    .io_cfg(OB1_io_cfg),
    .io_inputs_0(OB1_io_inputs_0),
    .io_outputs_0(OB1_io_outputs_0)
  );
  OB0 OB2 ( // @[TopModule.scala 220:48]
    .io_cfg(OB2_io_cfg),
    .io_inputs_0(OB2_io_inputs_0),
    .io_outputs_0(OB2_io_outputs_0)
  );
  OB0 OB3 ( // @[TopModule.scala 220:48]
    .io_cfg(OB3_io_cfg),
    .io_inputs_0(OB3_io_inputs_0),
    .io_outputs_0(OB3_io_outputs_0)
  );
  OB0 OB4 ( // @[TopModule.scala 220:48]
    .io_cfg(OB4_io_cfg),
    .io_inputs_0(OB4_io_inputs_0),
    .io_outputs_0(OB4_io_outputs_0)
  );
  OB0 OB5 ( // @[TopModule.scala 220:48]
    .io_cfg(OB5_io_cfg),
    .io_inputs_0(OB5_io_inputs_0),
    .io_outputs_0(OB5_io_outputs_0)
  );
  OB0 OB6 ( // @[TopModule.scala 220:48]
    .io_cfg(OB6_io_cfg),
    .io_inputs_0(OB6_io_inputs_0),
    .io_outputs_0(OB6_io_outputs_0)
  );
  OB0 OB7 ( // @[TopModule.scala 220:48]
    .io_cfg(OB7_io_cfg),
    .io_inputs_0(OB7_io_inputs_0),
    .io_outputs_0(OB7_io_outputs_0)
  );
  OB0 OB8 ( // @[TopModule.scala 220:48]
    .io_cfg(OB8_io_cfg),
    .io_inputs_0(OB8_io_inputs_0),
    .io_outputs_0(OB8_io_outputs_0)
  );
  OB0 OB9 ( // @[TopModule.scala 220:48]
    .io_cfg(OB9_io_cfg),
    .io_inputs_0(OB9_io_inputs_0),
    .io_outputs_0(OB9_io_outputs_0)
  );
  OB0 OB10 ( // @[TopModule.scala 220:48]
    .io_cfg(OB10_io_cfg),
    .io_inputs_0(OB10_io_inputs_0),
    .io_outputs_0(OB10_io_outputs_0)
  );
  OB0 OB11 ( // @[TopModule.scala 220:48]
    .io_cfg(OB11_io_cfg),
    .io_inputs_0(OB11_io_inputs_0),
    .io_outputs_0(OB11_io_outputs_0)
  );
  OB0 OB12 ( // @[TopModule.scala 220:48]
    .io_cfg(OB12_io_cfg),
    .io_inputs_0(OB12_io_inputs_0),
    .io_outputs_0(OB12_io_outputs_0)
  );
  OB0 OB13 ( // @[TopModule.scala 220:48]
    .io_cfg(OB13_io_cfg),
    .io_inputs_0(OB13_io_inputs_0),
    .io_outputs_0(OB13_io_outputs_0)
  );
  OB0 OB14 ( // @[TopModule.scala 220:48]
    .io_cfg(OB14_io_cfg),
    .io_inputs_0(OB14_io_inputs_0),
    .io_outputs_0(OB14_io_outputs_0)
  );
  OB0 OB15 ( // @[TopModule.scala 220:48]
    .io_cfg(OB15_io_cfg),
    .io_inputs_0(OB15_io_inputs_0),
    .io_outputs_0(OB15_io_outputs_0)
  );
  CfgMem_19 CfgMem ( // @[TopModule.scala 232:29]
    .clock(CfgMem_clock),
    .reset(CfgMem_reset),
    .io_cfgEn(CfgMem_io_cfgEn),
    .io_cfgData(CfgMem_io_cfgData),
    .io_cfgOut(CfgMem_io_cfgOut)
  );
  dpicCGRA dpicCGRA ( // @[TopModule.scala 292:27]
    .ins_0(dpicCGRA_ins_0),
    .ins_1(dpicCGRA_ins_1),
    .ins_2(dpicCGRA_ins_2),
    .ins_3(dpicCGRA_ins_3),
    .ins_4(dpicCGRA_ins_4),
    .ins_5(dpicCGRA_ins_5),
    .ins_6(dpicCGRA_ins_6),
    .ins_7(dpicCGRA_ins_7),
    .ins_8(dpicCGRA_ins_8),
    .ins_9(dpicCGRA_ins_9),
    .ins_10(dpicCGRA_ins_10),
    .ins_11(dpicCGRA_ins_11),
    .ins_12(dpicCGRA_ins_12),
    .ins_13(dpicCGRA_ins_13),
    .ins_14(dpicCGRA_ins_14),
    .ins_15(dpicCGRA_ins_15)
  );
  assign io_outputs_0 = OB0_io_outputs_0; // @[TopModule.scala 350:22]
  assign io_outputs_1 = OB1_io_outputs_0; // @[TopModule.scala 350:22]
  assign io_outputs_2 = OB2_io_outputs_0; // @[TopModule.scala 350:22]
  assign io_outputs_3 = OB3_io_outputs_0; // @[TopModule.scala 350:22]
  assign io_outputs_4 = OB4_io_outputs_0; // @[TopModule.scala 350:22]
  assign io_outputs_5 = OB5_io_outputs_0; // @[TopModule.scala 350:22]
  assign io_outputs_6 = OB6_io_outputs_0; // @[TopModule.scala 350:22]
  assign io_outputs_7 = OB7_io_outputs_0; // @[TopModule.scala 350:22]
  assign io_outputs_8 = OB8_io_outputs_0; // @[TopModule.scala 350:22]
  assign io_outputs_9 = OB9_io_outputs_0; // @[TopModule.scala 350:22]
  assign io_outputs_10 = OB10_io_outputs_0; // @[TopModule.scala 350:22]
  assign io_outputs_11 = OB11_io_outputs_0; // @[TopModule.scala 350:22]
  assign io_outputs_12 = OB12_io_outputs_0; // @[TopModule.scala 350:22]
  assign io_outputs_13 = OB13_io_outputs_0; // @[TopModule.scala 350:22]
  assign io_outputs_14 = OB14_io_outputs_0; // @[TopModule.scala 350:22]
  assign io_outputs_15 = OB15_io_outputs_0; // @[TopModule.scala 350:22]
  assign PE0_clock = clock;
  assign PE0_reset = reset;
  assign PE0_io_cfgEn = io_cfgEn & _T_1; // @[TopModule.scala 159:28]
  assign PE0_io_cfgData = io_cfgData; // @[TopModule.scala 161:30]
  assign PE0_io_inputs_0 = MatrixFC1_io_outputs_1; // @[TopModule.scala 350:22]
  assign PE0_io_inputs_1 = MatrixFC1_io_outputs_9; // @[TopModule.scala 350:22]
  assign PE1_clock = clock;
  assign PE1_reset = reset;
  assign PE1_io_cfgEn = io_cfgEn & _T_4; // @[TopModule.scala 159:28]
  assign PE1_io_cfgData = io_cfgData; // @[TopModule.scala 161:30]
  assign PE1_io_inputs_0 = MatrixFC1_io_outputs_2; // @[TopModule.scala 350:22]
  assign PE1_io_inputs_1 = MatrixFC1_io_outputs_10; // @[TopModule.scala 350:22]
  assign PE2_clock = clock;
  assign PE2_reset = reset;
  assign PE2_io_cfgEn = io_cfgEn & _T_7; // @[TopModule.scala 159:28]
  assign PE2_io_cfgData = io_cfgData; // @[TopModule.scala 161:30]
  assign PE2_io_inputs_0 = MatrixFC1_io_outputs_3; // @[TopModule.scala 350:22]
  assign PE2_io_inputs_1 = MatrixFC1_io_outputs_11; // @[TopModule.scala 350:22]
  assign PE3_clock = clock;
  assign PE3_reset = reset;
  assign PE3_io_cfgEn = io_cfgEn & _T_10; // @[TopModule.scala 159:28]
  assign PE3_io_cfgData = io_cfgData; // @[TopModule.scala 161:30]
  assign PE3_io_inputs_0 = MatrixFC1_io_outputs_4; // @[TopModule.scala 350:22]
  assign PE3_io_inputs_1 = MatrixFC1_io_outputs_12; // @[TopModule.scala 350:22]
  assign PE4_clock = clock;
  assign PE4_reset = reset;
  assign PE4_io_cfgEn = io_cfgEn & _T_13; // @[TopModule.scala 159:28]
  assign PE4_io_cfgData = io_cfgData; // @[TopModule.scala 161:30]
  assign PE4_io_inputs_0 = MatrixFC1_io_outputs_5; // @[TopModule.scala 350:22]
  assign PE4_io_inputs_1 = MatrixFC1_io_outputs_13; // @[TopModule.scala 350:22]
  assign PE5_clock = clock;
  assign PE5_reset = reset;
  assign PE5_io_cfgEn = io_cfgEn & _T_16; // @[TopModule.scala 159:28]
  assign PE5_io_cfgData = io_cfgData; // @[TopModule.scala 161:30]
  assign PE5_io_inputs_0 = MatrixFC1_io_outputs_6; // @[TopModule.scala 350:22]
  assign PE5_io_inputs_1 = MatrixFC1_io_outputs_14; // @[TopModule.scala 350:22]
  assign PE6_clock = clock;
  assign PE6_reset = reset;
  assign PE6_io_cfgEn = io_cfgEn & _T_19; // @[TopModule.scala 159:28]
  assign PE6_io_cfgData = io_cfgData; // @[TopModule.scala 161:30]
  assign PE6_io_inputs_0 = MatrixFC1_io_outputs_7; // @[TopModule.scala 350:22]
  assign PE6_io_inputs_1 = MatrixFC1_io_outputs_15; // @[TopModule.scala 350:22]
  assign PE7_clock = clock;
  assign PE7_reset = reset;
  assign PE7_io_cfgEn = io_cfgEn & _T_22; // @[TopModule.scala 159:28]
  assign PE7_io_cfgData = io_cfgData; // @[TopModule.scala 161:30]
  assign PE7_io_inputs_0 = MatrixFC1_io_outputs_8; // @[TopModule.scala 350:22]
  assign PE7_io_inputs_1 = MatrixFC1_io_outputs_16; // @[TopModule.scala 350:22]
  assign PE8_clock = clock;
  assign PE8_reset = reset;
  assign PE8_io_cfgEn = io_cfgEn & _T_25; // @[TopModule.scala 159:28]
  assign PE8_io_cfgData = io_cfgData; // @[TopModule.scala 161:30]
  assign PE8_io_inputs_0 = MatrixFC0_io_outputs_1; // @[TopModule.scala 350:22]
  assign PE8_io_inputs_1 = MatrixFC0_io_outputs_9; // @[TopModule.scala 350:22]
  assign dpicDebug_in = PE8_io_outputs_0; // @[TopModule.scala 166:27]
  assign PE9_clock = clock;
  assign PE9_reset = reset;
  assign PE9_io_cfgEn = io_cfgEn & _T_28; // @[TopModule.scala 159:28]
  assign PE9_io_cfgData = io_cfgData; // @[TopModule.scala 161:30]
  assign PE9_io_inputs_0 = MatrixFC0_io_outputs_2; // @[TopModule.scala 350:22]
  assign PE9_io_inputs_1 = MatrixFC0_io_outputs_10; // @[TopModule.scala 350:22]
  assign PE10_clock = clock;
  assign PE10_reset = reset;
  assign PE10_io_cfgEn = io_cfgEn & _T_31; // @[TopModule.scala 159:28]
  assign PE10_io_cfgData = io_cfgData; // @[TopModule.scala 161:30]
  assign PE10_io_inputs_0 = MatrixFC0_io_outputs_3; // @[TopModule.scala 350:22]
  assign PE10_io_inputs_1 = MatrixFC0_io_outputs_11; // @[TopModule.scala 350:22]
  assign PE11_clock = clock;
  assign PE11_reset = reset;
  assign PE11_io_cfgEn = io_cfgEn & _T_34; // @[TopModule.scala 159:28]
  assign PE11_io_cfgData = io_cfgData; // @[TopModule.scala 161:30]
  assign PE11_io_inputs_0 = MatrixFC0_io_outputs_4; // @[TopModule.scala 350:22]
  assign PE11_io_inputs_1 = MatrixFC0_io_outputs_12; // @[TopModule.scala 350:22]
  assign PE12_clock = clock;
  assign PE12_reset = reset;
  assign PE12_io_cfgEn = io_cfgEn & _T_37; // @[TopModule.scala 159:28]
  assign PE12_io_cfgData = io_cfgData; // @[TopModule.scala 161:30]
  assign PE12_io_inputs_0 = MatrixFC0_io_outputs_5; // @[TopModule.scala 350:22]
  assign PE12_io_inputs_1 = MatrixFC0_io_outputs_13; // @[TopModule.scala 350:22]
  assign PE13_clock = clock;
  assign PE13_reset = reset;
  assign PE13_io_cfgEn = io_cfgEn & _T_40; // @[TopModule.scala 159:28]
  assign PE13_io_cfgData = io_cfgData; // @[TopModule.scala 161:30]
  assign PE13_io_inputs_0 = MatrixFC0_io_outputs_6; // @[TopModule.scala 350:22]
  assign PE13_io_inputs_1 = MatrixFC0_io_outputs_14; // @[TopModule.scala 350:22]
  assign PE14_clock = clock;
  assign PE14_reset = reset;
  assign PE14_io_cfgEn = io_cfgEn & _T_43; // @[TopModule.scala 159:28]
  assign PE14_io_cfgData = io_cfgData; // @[TopModule.scala 161:30]
  assign PE14_io_inputs_0 = MatrixFC0_io_outputs_7; // @[TopModule.scala 350:22]
  assign PE14_io_inputs_1 = MatrixFC0_io_outputs_15; // @[TopModule.scala 350:22]
  assign PE15_clock = clock;
  assign PE15_reset = reset;
  assign PE15_io_cfgEn = io_cfgEn & _T_46; // @[TopModule.scala 159:28]
  assign PE15_io_cfgData = io_cfgData; // @[TopModule.scala 161:30]
  assign PE15_io_inputs_0 = MatrixFC0_io_outputs_8; // @[TopModule.scala 350:22]
  assign PE15_io_inputs_1 = MatrixFC0_io_outputs_16; // @[TopModule.scala 350:22]
  assign MatrixFC0_clock = clock;
  assign MatrixFC0_reset = reset;
  assign MatrixFC0_io_cfgEn = io_cfgEn & _T_49; // @[TopModule.scala 159:28]
  assign MatrixFC0_io_cfgAddr = io_cfgAddr[3:0]; // @[TopModule.scala 160:30]
  assign MatrixFC0_io_cfgData = io_cfgData; // @[TopModule.scala 161:30]
  assign MatrixFC0_io_inputs_0 = MatrixFC1_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC0_io_inputs_1 = PE0_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC0_io_inputs_2 = PE1_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC0_io_inputs_3 = PE2_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC0_io_inputs_4 = PE3_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC0_io_inputs_5 = PE4_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC0_io_inputs_6 = PE5_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC0_io_inputs_7 = PE6_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC0_io_inputs_8 = PE7_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC0_io_inputs_9 = PE8_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC0_io_inputs_10 = PE9_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC0_io_inputs_11 = PE10_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC0_io_inputs_12 = PE11_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC0_io_inputs_13 = PE12_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC0_io_inputs_14 = PE13_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC0_io_inputs_15 = PE14_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC0_io_inputs_16 = PE15_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_clock = clock;
  assign MatrixFC1_reset = reset;
  assign MatrixFC1_io_cfgEn = io_cfgEn & _T_52; // @[TopModule.scala 159:28]
  assign MatrixFC1_io_cfgAddr = io_cfgAddr[3:0]; // @[TopModule.scala 160:30]
  assign MatrixFC1_io_cfgData = io_cfgData; // @[TopModule.scala 161:30]
  assign MatrixFC1_io_inputs_0 = IB0_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_1 = IB1_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_2 = IB2_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_3 = IB3_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_4 = IB4_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_5 = IB5_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_6 = IB6_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_7 = IB7_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_8 = IB8_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_9 = IB9_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_10 = IB10_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_11 = IB11_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_12 = IB12_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_13 = IB13_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_14 = IB14_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_15 = IB15_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_16 = PE0_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_17 = PE1_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_18 = PE2_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_19 = PE3_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_20 = PE4_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_21 = PE5_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_22 = PE6_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC1_io_inputs_23 = PE7_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC2_clock = clock;
  assign MatrixFC2_reset = reset;
  assign MatrixFC2_io_cfgEn = io_cfgEn & _T_55; // @[TopModule.scala 159:28]
  assign MatrixFC2_io_cfgAddr = io_cfgAddr[3:0]; // @[TopModule.scala 160:30]
  assign MatrixFC2_io_cfgData = io_cfgData; // @[TopModule.scala 161:30]
  assign MatrixFC2_io_inputs_0 = MatrixFC0_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC2_io_inputs_1 = PE8_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC2_io_inputs_2 = PE9_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC2_io_inputs_3 = PE10_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC2_io_inputs_4 = PE11_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC2_io_inputs_5 = PE12_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC2_io_inputs_6 = PE13_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC2_io_inputs_7 = PE14_io_outputs_0; // @[TopModule.scala 350:22]
  assign MatrixFC2_io_inputs_8 = PE15_io_outputs_0; // @[TopModule.scala 350:22]
  assign IB0_io_inputs_0 = io_inputs_0; // @[TopModule.scala 350:22]
  assign IB1_io_inputs_0 = io_inputs_1; // @[TopModule.scala 350:22]
  assign IB2_io_inputs_0 = io_inputs_2; // @[TopModule.scala 350:22]
  assign IB3_io_inputs_0 = io_inputs_3; // @[TopModule.scala 350:22]
  assign IB4_io_inputs_0 = io_inputs_4; // @[TopModule.scala 350:22]
  assign IB5_io_inputs_0 = io_inputs_5; // @[TopModule.scala 350:22]
  assign IB6_io_inputs_0 = io_inputs_6; // @[TopModule.scala 350:22]
  assign IB7_io_inputs_0 = io_inputs_7; // @[TopModule.scala 350:22]
  assign IB8_io_inputs_0 = io_inputs_8; // @[TopModule.scala 350:22]
  assign IB9_io_inputs_0 = io_inputs_9; // @[TopModule.scala 350:22]
  assign IB10_io_inputs_0 = io_inputs_10; // @[TopModule.scala 350:22]
  assign IB11_io_inputs_0 = io_inputs_11; // @[TopModule.scala 350:22]
  assign IB12_io_inputs_0 = io_inputs_12; // @[TopModule.scala 350:22]
  assign IB13_io_inputs_0 = io_inputs_13; // @[TopModule.scala 350:22]
  assign IB14_io_inputs_0 = io_inputs_14; // @[TopModule.scala 350:22]
  assign IB15_io_inputs_0 = io_inputs_15; // @[TopModule.scala 350:22]
  assign OB0_io_cfg = CfgMem_io_cfgOut[0]; // @[TopModule.scala 263:80]
  assign OB0_io_inputs_0 = MatrixFC2_io_outputs_0; // @[TopModule.scala 350:22]
  assign OB1_io_cfg = CfgMem_io_cfgOut[1]; // @[TopModule.scala 263:80]
  assign OB1_io_inputs_0 = MatrixFC2_io_outputs_1; // @[TopModule.scala 350:22]
  assign OB2_io_cfg = CfgMem_io_cfgOut[2]; // @[TopModule.scala 263:80]
  assign OB2_io_inputs_0 = MatrixFC2_io_outputs_2; // @[TopModule.scala 350:22]
  assign OB3_io_cfg = CfgMem_io_cfgOut[3]; // @[TopModule.scala 263:80]
  assign OB3_io_inputs_0 = MatrixFC2_io_outputs_3; // @[TopModule.scala 350:22]
  assign OB4_io_cfg = CfgMem_io_cfgOut[4]; // @[TopModule.scala 263:80]
  assign OB4_io_inputs_0 = MatrixFC2_io_outputs_4; // @[TopModule.scala 350:22]
  assign OB5_io_cfg = CfgMem_io_cfgOut[5]; // @[TopModule.scala 263:80]
  assign OB5_io_inputs_0 = MatrixFC2_io_outputs_5; // @[TopModule.scala 350:22]
  assign OB6_io_cfg = CfgMem_io_cfgOut[6]; // @[TopModule.scala 263:80]
  assign OB6_io_inputs_0 = MatrixFC2_io_outputs_6; // @[TopModule.scala 350:22]
  assign OB7_io_cfg = CfgMem_io_cfgOut[7]; // @[TopModule.scala 263:80]
  assign OB7_io_inputs_0 = MatrixFC2_io_outputs_7; // @[TopModule.scala 350:22]
  assign OB8_io_cfg = CfgMem_io_cfgOut[8]; // @[TopModule.scala 263:80]
  assign OB8_io_inputs_0 = MatrixFC2_io_outputs_8; // @[TopModule.scala 350:22]
  assign OB9_io_cfg = CfgMem_io_cfgOut[9]; // @[TopModule.scala 263:80]
  assign OB9_io_inputs_0 = MatrixFC2_io_outputs_9; // @[TopModule.scala 350:22]
  assign OB10_io_cfg = CfgMem_io_cfgOut[10]; // @[TopModule.scala 263:80]
  assign OB10_io_inputs_0 = MatrixFC2_io_outputs_10; // @[TopModule.scala 350:22]
  assign OB11_io_cfg = CfgMem_io_cfgOut[11]; // @[TopModule.scala 263:80]
  assign OB11_io_inputs_0 = MatrixFC2_io_outputs_11; // @[TopModule.scala 350:22]
  assign OB12_io_cfg = CfgMem_io_cfgOut[12]; // @[TopModule.scala 263:80]
  assign OB12_io_inputs_0 = MatrixFC2_io_outputs_12; // @[TopModule.scala 350:22]
  assign OB13_io_cfg = CfgMem_io_cfgOut[13]; // @[TopModule.scala 263:80]
  assign OB13_io_inputs_0 = MatrixFC2_io_outputs_13; // @[TopModule.scala 350:22]
  assign OB14_io_cfg = CfgMem_io_cfgOut[14]; // @[TopModule.scala 263:80]
  assign OB14_io_inputs_0 = MatrixFC2_io_outputs_14; // @[TopModule.scala 350:22]
  assign OB15_io_cfg = CfgMem_io_cfgOut[15]; // @[TopModule.scala 263:80]
  assign OB15_io_inputs_0 = MatrixFC2_io_outputs_15; // @[TopModule.scala 350:22]
  assign CfgMem_clock = clock;
  assign CfgMem_reset = reset;
  assign CfgMem_io_cfgEn = io_cfgEn & _T_58; // @[TopModule.scala 241:34]
  assign CfgMem_io_cfgData = io_cfgData; // @[TopModule.scala 248:28]
  assign dpicCGRA_ins_0 = io_inputs_0; // @[TopModule.scala 297:31]
  assign dpicCGRA_ins_1 = io_inputs_1; // @[TopModule.scala 297:31]
  assign dpicCGRA_ins_2 = io_inputs_2; // @[TopModule.scala 297:31]
  assign dpicCGRA_ins_3 = io_inputs_3; // @[TopModule.scala 297:31]
  assign dpicCGRA_ins_4 = io_inputs_4; // @[TopModule.scala 297:31]
  assign dpicCGRA_ins_5 = io_inputs_5; // @[TopModule.scala 297:31]
  assign dpicCGRA_ins_6 = io_inputs_6; // @[TopModule.scala 297:31]
  assign dpicCGRA_ins_7 = io_inputs_7; // @[TopModule.scala 297:31]
  assign dpicCGRA_ins_8 = io_inputs_8; // @[TopModule.scala 297:31]
  assign dpicCGRA_ins_9 = io_inputs_9; // @[TopModule.scala 297:31]
  assign dpicCGRA_ins_10 = io_inputs_10; // @[TopModule.scala 297:31]
  assign dpicCGRA_ins_11 = io_inputs_11; // @[TopModule.scala 297:31]
  assign dpicCGRA_ins_12 = io_inputs_12; // @[TopModule.scala 297:31]
  assign dpicCGRA_ins_13 = io_inputs_13; // @[TopModule.scala 297:31]
  assign dpicCGRA_ins_14 = io_inputs_14; // @[TopModule.scala 297:31]
  assign dpicCGRA_ins_15 = io_inputs_15; // @[TopModule.scala 297:31]
endmodule
module CGRAFullMask(
  input          clock,
  input          reset,
  input          io_CGRAIO_valid,
  output         io_CGRAIO_ready,
  output [63:0]  io_CGRAIO_data_read,
  input  [63:0]  io_CGRAIO_data_write,
  input          io_CGRAIO_wen,
  input  [31:0]  io_CGRAIO_addr,
  output [32:0]  io_outputs_0,
  output [32:0]  io_outputs_1,
  output [32:0]  io_outputs_2,
  output [32:0]  io_outputs_3,
  output [32:0]  io_outputs_4,
  output [32:0]  io_outputs_5,
  output [32:0]  io_outputs_6,
  output [32:0]  io_outputs_7,
  output [32:0]  io_outputs_8,
  output [32:0]  io_outputs_9,
  output [32:0]  io_outputs_10,
  output [32:0]  io_outputs_11,
  output [32:0]  io_outputs_12,
  output [32:0]  io_outputs_13,
  output [32:0]  io_outputs_14,
  output [32:0]  io_outputs_15,
  input          _T_100_0,
  input  [191:0] dmaCtrl
);
  wire  outQueue_0_clock; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_0_reset; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_0_io_enq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_0_io_enq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_0_io_enq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_0_io_deq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_0_io_deq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_0_io_deq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_1_clock; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_1_reset; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_1_io_enq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_1_io_enq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_1_io_enq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_1_io_deq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_1_io_deq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_1_io_deq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_2_clock; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_2_reset; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_2_io_enq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_2_io_enq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_2_io_enq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_2_io_deq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_2_io_deq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_2_io_deq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_3_clock; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_3_reset; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_3_io_enq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_3_io_enq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_3_io_enq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_3_io_deq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_3_io_deq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_3_io_deq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_4_clock; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_4_reset; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_4_io_enq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_4_io_enq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_4_io_enq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_4_io_deq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_4_io_deq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_4_io_deq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_5_clock; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_5_reset; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_5_io_enq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_5_io_enq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_5_io_enq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_5_io_deq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_5_io_deq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_5_io_deq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_6_clock; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_6_reset; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_6_io_enq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_6_io_enq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_6_io_enq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_6_io_deq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_6_io_deq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_6_io_deq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_7_clock; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_7_reset; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_7_io_enq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_7_io_enq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_7_io_enq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_7_io_deq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_7_io_deq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_7_io_deq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_8_clock; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_8_reset; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_8_io_enq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_8_io_enq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_8_io_enq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_8_io_deq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_8_io_deq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_8_io_deq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_9_clock; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_9_reset; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_9_io_enq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_9_io_enq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_9_io_enq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_9_io_deq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_9_io_deq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_9_io_deq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_10_clock; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_10_reset; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_10_io_enq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_10_io_enq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_10_io_enq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_10_io_deq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_10_io_deq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_10_io_deq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_11_clock; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_11_reset; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_11_io_enq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_11_io_enq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_11_io_enq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_11_io_deq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_11_io_deq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_11_io_deq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_12_clock; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_12_reset; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_12_io_enq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_12_io_enq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_12_io_enq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_12_io_deq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_12_io_deq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_12_io_deq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_13_clock; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_13_reset; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_13_io_enq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_13_io_enq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_13_io_enq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_13_io_deq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_13_io_deq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_13_io_deq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_14_clock; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_14_reset; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_14_io_enq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_14_io_enq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_14_io_enq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_14_io_deq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_14_io_deq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_14_io_deq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_15_clock; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_15_reset; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_15_io_enq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_15_io_enq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_15_io_enq_bits; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_15_io_deq_ready; // @[CGRAFullMask.scala 16:52]
  wire  outQueue_15_io_deq_valid; // @[CGRAFullMask.scala 16:52]
  wire [31:0] outQueue_15_io_deq_bits; // @[CGRAFullMask.scala 16:52]
  wire  synInInst_clock; // @[CGRAFullMask.scala 19:25]
  wire  synInInst_reset; // @[CGRAFullMask.scala 19:25]
  wire  synInInst_io_valid; // @[CGRAFullMask.scala 19:25]
  wire  synInInst_io_ready; // @[CGRAFullMask.scala 19:25]
  wire [63:0] synInInst_io_dataIn; // @[CGRAFullMask.scala 19:25]
  wire [32:0] synInInst_io_dataOut_0; // @[CGRAFullMask.scala 19:25]
  wire [32:0] synInInst_io_dataOut_1; // @[CGRAFullMask.scala 19:25]
  wire [32:0] synInInst_io_dataOut_2; // @[CGRAFullMask.scala 19:25]
  wire [32:0] synInInst_io_dataOut_3; // @[CGRAFullMask.scala 19:25]
  wire [32:0] synInInst_io_dataOut_4; // @[CGRAFullMask.scala 19:25]
  wire [32:0] synInInst_io_dataOut_5; // @[CGRAFullMask.scala 19:25]
  wire [32:0] synInInst_io_dataOut_6; // @[CGRAFullMask.scala 19:25]
  wire [32:0] synInInst_io_dataOut_7; // @[CGRAFullMask.scala 19:25]
  wire [32:0] synInInst_io_dataOut_8; // @[CGRAFullMask.scala 19:25]
  wire [32:0] synInInst_io_dataOut_9; // @[CGRAFullMask.scala 19:25]
  wire [32:0] synInInst_io_dataOut_10; // @[CGRAFullMask.scala 19:25]
  wire [32:0] synInInst_io_dataOut_11; // @[CGRAFullMask.scala 19:25]
  wire [32:0] synInInst_io_dataOut_12; // @[CGRAFullMask.scala 19:25]
  wire [32:0] synInInst_io_dataOut_13; // @[CGRAFullMask.scala 19:25]
  wire [32:0] synInInst_io_dataOut_14; // @[CGRAFullMask.scala 19:25]
  wire [32:0] synInInst_io_dataOut_15; // @[CGRAFullMask.scala 19:25]
  wire  synInInst_io_delayen; // @[CGRAFullMask.scala 19:25]
  wire [63:0] synInInst_io_delayCycle; // @[CGRAFullMask.scala 19:25]
  wire  synInInst_dmaEnWR_0; // @[CGRAFullMask.scala 19:25]
  wire [191:0] synInInst_dmaCtrl_0; // @[CGRAFullMask.scala 19:25]
  wire  cgraInst_clock; // @[CGRAFullMask.scala 23:35]
  wire  cgraInst_reset; // @[CGRAFullMask.scala 23:35]
  wire  cgraInst_io_cfgEn; // @[CGRAFullMask.scala 23:35]
  wire [8:0] cgraInst_io_cfgAddr; // @[CGRAFullMask.scala 23:35]
  wire [31:0] cgraInst_io_cfgData; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_inputs_0; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_inputs_1; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_inputs_2; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_inputs_3; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_inputs_4; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_inputs_5; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_inputs_6; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_inputs_7; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_inputs_8; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_inputs_9; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_inputs_10; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_inputs_11; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_inputs_12; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_inputs_13; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_inputs_14; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_inputs_15; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_outputs_0; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_outputs_1; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_outputs_2; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_outputs_3; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_outputs_4; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_outputs_5; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_outputs_6; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_outputs_7; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_outputs_8; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_outputs_9; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_outputs_10; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_outputs_11; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_outputs_12; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_outputs_13; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_outputs_14; // @[CGRAFullMask.scala 23:35]
  wire [32:0] cgraInst_io_outputs_15; // @[CGRAFullMask.scala 23:35]
  wire  _T_32 = io_CGRAIO_addr >= 32'h2010000; // @[CGRAFullMask.scala 33:32]
  wire  _T_35 = io_CGRAIO_addr <= 32'h2010040; // @[CGRAFullMask.scala 33:67]
  wire  addrIsW = _T_32 & _T_35; // @[CGRAFullMask.scala 33:49]
  wire  oneHList2_0 = 32'h2010040 == io_CGRAIO_addr; // @[CGRAFullMask.scala 39:46]
  wire  oneHList2_1 = 32'h2010044 == io_CGRAIO_addr; // @[CGRAFullMask.scala 39:46]
  wire  oneHList2_2 = 32'h2010048 == io_CGRAIO_addr; // @[CGRAFullMask.scala 39:46]
  wire  oneHList2_3 = 32'h201004c == io_CGRAIO_addr; // @[CGRAFullMask.scala 39:46]
  wire  oneHList2_4 = 32'h2010050 == io_CGRAIO_addr; // @[CGRAFullMask.scala 39:46]
  wire  oneHList2_5 = 32'h2010054 == io_CGRAIO_addr; // @[CGRAFullMask.scala 39:46]
  wire  oneHList2_6 = 32'h2010058 == io_CGRAIO_addr; // @[CGRAFullMask.scala 39:46]
  wire  oneHList2_7 = 32'h201005c == io_CGRAIO_addr; // @[CGRAFullMask.scala 39:46]
  wire  oneHList2_8 = 32'h2010060 == io_CGRAIO_addr; // @[CGRAFullMask.scala 39:46]
  wire  oneHList2_9 = 32'h2010064 == io_CGRAIO_addr; // @[CGRAFullMask.scala 39:46]
  wire  oneHList2_10 = 32'h2010068 == io_CGRAIO_addr; // @[CGRAFullMask.scala 39:46]
  wire  oneHList2_11 = 32'h201006c == io_CGRAIO_addr; // @[CGRAFullMask.scala 39:46]
  wire  oneHList2_12 = 32'h2010070 == io_CGRAIO_addr; // @[CGRAFullMask.scala 39:46]
  wire  oneHList2_13 = 32'h2010074 == io_CGRAIO_addr; // @[CGRAFullMask.scala 39:46]
  wire  oneHList2_14 = 32'h2010078 == io_CGRAIO_addr; // @[CGRAFullMask.scala 39:46]
  wire  oneHList2_15 = 32'h201007c == io_CGRAIO_addr; // @[CGRAFullMask.scala 39:46]
  wire  oneHot_17 = 32'h2010080 == io_CGRAIO_addr; // @[CGRAFullMask.scala 43:116]
  wire  oneHot_18 = 32'h2010088 == io_CGRAIO_addr; // @[CGRAFullMask.scala 44:83]
  wire [9:0] _T_88 = {addrIsW,oneHList2_0,oneHList2_1,oneHList2_2,oneHList2_3,oneHList2_4,oneHList2_5,oneHList2_6,oneHList2_7,oneHList2_8}; // @[Cat.scala 29:58]
  wire [18:0] _T_89 = {_T_88,oneHList2_9,oneHList2_10,oneHList2_11,oneHList2_12,oneHList2_13,oneHList2_14,oneHList2_15,oneHot_17,oneHot_18}; // @[Cat.scala 29:58]
  wire [9:0] _T_106 = {synInInst_io_ready,outQueue_0_io_deq_valid,outQueue_1_io_deq_valid,outQueue_2_io_deq_valid,outQueue_3_io_deq_valid,outQueue_4_io_deq_valid,outQueue_5_io_deq_valid,outQueue_6_io_deq_valid,outQueue_7_io_deq_valid,outQueue_8_io_deq_valid}; // @[Cat.scala 29:58]
  wire [18:0] _T_107 = {_T_106,outQueue_9_io_deq_valid,outQueue_10_io_deq_valid,outQueue_11_io_deq_valid,outQueue_12_io_deq_valid,outQueue_13_io_deq_valid,outQueue_14_io_deq_valid,outQueue_15_io_deq_valid,2'h3}; // @[Cat.scala 29:58]
  wire  _T_108 = addrIsW & synInInst_io_ready; // @[Mux.scala 27:72]
  wire  _T_109 = oneHList2_0 & outQueue_0_io_deq_valid; // @[Mux.scala 27:72]
  wire  _T_110 = oneHList2_1 & outQueue_1_io_deq_valid; // @[Mux.scala 27:72]
  wire  _T_111 = oneHList2_2 & outQueue_2_io_deq_valid; // @[Mux.scala 27:72]
  wire  _T_112 = oneHList2_3 & outQueue_3_io_deq_valid; // @[Mux.scala 27:72]
  wire  _T_113 = oneHList2_4 & outQueue_4_io_deq_valid; // @[Mux.scala 27:72]
  wire  _T_114 = oneHList2_5 & outQueue_5_io_deq_valid; // @[Mux.scala 27:72]
  wire  _T_115 = oneHList2_6 & outQueue_6_io_deq_valid; // @[Mux.scala 27:72]
  wire  _T_116 = oneHList2_7 & outQueue_7_io_deq_valid; // @[Mux.scala 27:72]
  wire  _T_117 = oneHList2_8 & outQueue_8_io_deq_valid; // @[Mux.scala 27:72]
  wire  _T_118 = oneHList2_9 & outQueue_9_io_deq_valid; // @[Mux.scala 27:72]
  wire  _T_119 = oneHList2_10 & outQueue_10_io_deq_valid; // @[Mux.scala 27:72]
  wire  _T_120 = oneHList2_11 & outQueue_11_io_deq_valid; // @[Mux.scala 27:72]
  wire  _T_121 = oneHList2_12 & outQueue_12_io_deq_valid; // @[Mux.scala 27:72]
  wire  _T_122 = oneHList2_13 & outQueue_13_io_deq_valid; // @[Mux.scala 27:72]
  wire  _T_123 = oneHList2_14 & outQueue_14_io_deq_valid; // @[Mux.scala 27:72]
  wire  _T_124 = oneHList2_15 & outQueue_15_io_deq_valid; // @[Mux.scala 27:72]
  wire  _T_127 = _T_108 | _T_109; // @[Mux.scala 27:72]
  wire  _T_128 = _T_127 | _T_110; // @[Mux.scala 27:72]
  wire  _T_129 = _T_128 | _T_111; // @[Mux.scala 27:72]
  wire  _T_130 = _T_129 | _T_112; // @[Mux.scala 27:72]
  wire  _T_131 = _T_130 | _T_113; // @[Mux.scala 27:72]
  wire  _T_132 = _T_131 | _T_114; // @[Mux.scala 27:72]
  wire  _T_133 = _T_132 | _T_115; // @[Mux.scala 27:72]
  wire  _T_134 = _T_133 | _T_116; // @[Mux.scala 27:72]
  wire  _T_135 = _T_134 | _T_117; // @[Mux.scala 27:72]
  wire  _T_136 = _T_135 | _T_118; // @[Mux.scala 27:72]
  wire  _T_137 = _T_136 | _T_119; // @[Mux.scala 27:72]
  wire  _T_138 = _T_137 | _T_120; // @[Mux.scala 27:72]
  wire  _T_139 = _T_138 | _T_121; // @[Mux.scala 27:72]
  wire  _T_140 = _T_139 | _T_122; // @[Mux.scala 27:72]
  wire  _T_141 = _T_140 | _T_123; // @[Mux.scala 27:72]
  wire  _T_142 = _T_141 | _T_124; // @[Mux.scala 27:72]
  wire  _T_143 = _T_142 | oneHot_17; // @[Mux.scala 27:72]
  wire  _T_146 = io_CGRAIO_valid & io_CGRAIO_wen; // @[CGRAFullMask.scala 65:41]
  wire  _T_150 = io_CGRAIO_addr == 32'h2010040; // @[CGRAFullMask.scala 67:53]
  wire  _T_154 = io_CGRAIO_addr == 32'h2010044; // @[CGRAFullMask.scala 67:53]
  wire  _T_158 = io_CGRAIO_addr == 32'h2010048; // @[CGRAFullMask.scala 67:53]
  wire  _T_162 = io_CGRAIO_addr == 32'h201004c; // @[CGRAFullMask.scala 67:53]
  wire  _T_166 = io_CGRAIO_addr == 32'h2010050; // @[CGRAFullMask.scala 67:53]
  wire  _T_170 = io_CGRAIO_addr == 32'h2010054; // @[CGRAFullMask.scala 67:53]
  wire  _T_174 = io_CGRAIO_addr == 32'h2010058; // @[CGRAFullMask.scala 67:53]
  wire  _T_178 = io_CGRAIO_addr == 32'h201005c; // @[CGRAFullMask.scala 67:53]
  wire  _T_182 = io_CGRAIO_addr == 32'h2010060; // @[CGRAFullMask.scala 67:53]
  wire  _T_186 = io_CGRAIO_addr == 32'h2010064; // @[CGRAFullMask.scala 67:53]
  wire  _T_190 = io_CGRAIO_addr == 32'h2010068; // @[CGRAFullMask.scala 67:53]
  wire  _T_194 = io_CGRAIO_addr == 32'h201006c; // @[CGRAFullMask.scala 67:53]
  wire  _T_198 = io_CGRAIO_addr == 32'h2010070; // @[CGRAFullMask.scala 67:53]
  wire  _T_202 = io_CGRAIO_addr == 32'h2010074; // @[CGRAFullMask.scala 67:53]
  wire  _T_206 = io_CGRAIO_addr == 32'h2010078; // @[CGRAFullMask.scala 67:53]
  wire  _T_210 = io_CGRAIO_addr == 32'h201007c; // @[CGRAFullMask.scala 67:53]
  wire  _T_214 = io_CGRAIO_addr == 32'h2010080; // @[CGRAFullMask.scala 69:39]
  wire  _T_218 = io_CGRAIO_addr == 32'h2010088; // @[CGRAFullMask.scala 70:42]
  wire [31:0] _T_222 = oneHList2_0 ? outQueue_0_io_deq_bits : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_223 = oneHList2_1 ? outQueue_1_io_deq_bits : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_224 = oneHList2_2 ? outQueue_2_io_deq_bits : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_225 = oneHList2_3 ? outQueue_3_io_deq_bits : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_226 = oneHList2_4 ? outQueue_4_io_deq_bits : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_227 = oneHList2_5 ? outQueue_5_io_deq_bits : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_228 = oneHList2_6 ? outQueue_6_io_deq_bits : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_229 = oneHList2_7 ? outQueue_7_io_deq_bits : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_230 = oneHList2_8 ? outQueue_8_io_deq_bits : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_231 = oneHList2_9 ? outQueue_9_io_deq_bits : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_232 = oneHList2_10 ? outQueue_10_io_deq_bits : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_233 = oneHList2_11 ? outQueue_11_io_deq_bits : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_234 = oneHList2_12 ? outQueue_12_io_deq_bits : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_235 = oneHList2_13 ? outQueue_13_io_deq_bits : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_236 = oneHList2_14 ? outQueue_14_io_deq_bits : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_237 = oneHList2_15 ? outQueue_15_io_deq_bits : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_238 = _T_222 | _T_223; // @[Mux.scala 27:72]
  wire [31:0] _T_239 = _T_238 | _T_224; // @[Mux.scala 27:72]
  wire [31:0] _T_240 = _T_239 | _T_225; // @[Mux.scala 27:72]
  wire [31:0] _T_241 = _T_240 | _T_226; // @[Mux.scala 27:72]
  wire [31:0] _T_242 = _T_241 | _T_227; // @[Mux.scala 27:72]
  wire [31:0] _T_243 = _T_242 | _T_228; // @[Mux.scala 27:72]
  wire [31:0] _T_244 = _T_243 | _T_229; // @[Mux.scala 27:72]
  wire [31:0] _T_245 = _T_244 | _T_230; // @[Mux.scala 27:72]
  wire [31:0] _T_246 = _T_245 | _T_231; // @[Mux.scala 27:72]
  wire [31:0] _T_247 = _T_246 | _T_232; // @[Mux.scala 27:72]
  wire [31:0] _T_248 = _T_247 | _T_233; // @[Mux.scala 27:72]
  wire [31:0] _T_249 = _T_248 | _T_234; // @[Mux.scala 27:72]
  wire [31:0] _T_250 = _T_249 | _T_235; // @[Mux.scala 27:72]
  wire [31:0] _T_251 = _T_250 | _T_236; // @[Mux.scala 27:72]
  wire [31:0] _T_252 = _T_251 | _T_237; // @[Mux.scala 27:72]
  wire [18:0] oneHotWire = _T_89; // @[CGRAFullMask.scala 41:34 CGRAFullMask.scala 51:14]
  wire [18:0] outReadyList = _T_107; // @[CGRAFullMask.scala 42:35 CGRAFullMask.scala 52:16]
  Queue outQueue_0 ( // @[CGRAFullMask.scala 16:52]
    .clock(outQueue_0_clock),
    .reset(outQueue_0_reset),
    .io_enq_ready(outQueue_0_io_enq_ready),
    .io_enq_valid(outQueue_0_io_enq_valid),
    .io_enq_bits(outQueue_0_io_enq_bits),
    .io_deq_ready(outQueue_0_io_deq_ready),
    .io_deq_valid(outQueue_0_io_deq_valid),
    .io_deq_bits(outQueue_0_io_deq_bits)
  );
  Queue outQueue_1 ( // @[CGRAFullMask.scala 16:52]
    .clock(outQueue_1_clock),
    .reset(outQueue_1_reset),
    .io_enq_ready(outQueue_1_io_enq_ready),
    .io_enq_valid(outQueue_1_io_enq_valid),
    .io_enq_bits(outQueue_1_io_enq_bits),
    .io_deq_ready(outQueue_1_io_deq_ready),
    .io_deq_valid(outQueue_1_io_deq_valid),
    .io_deq_bits(outQueue_1_io_deq_bits)
  );
  Queue outQueue_2 ( // @[CGRAFullMask.scala 16:52]
    .clock(outQueue_2_clock),
    .reset(outQueue_2_reset),
    .io_enq_ready(outQueue_2_io_enq_ready),
    .io_enq_valid(outQueue_2_io_enq_valid),
    .io_enq_bits(outQueue_2_io_enq_bits),
    .io_deq_ready(outQueue_2_io_deq_ready),
    .io_deq_valid(outQueue_2_io_deq_valid),
    .io_deq_bits(outQueue_2_io_deq_bits)
  );
  Queue outQueue_3 ( // @[CGRAFullMask.scala 16:52]
    .clock(outQueue_3_clock),
    .reset(outQueue_3_reset),
    .io_enq_ready(outQueue_3_io_enq_ready),
    .io_enq_valid(outQueue_3_io_enq_valid),
    .io_enq_bits(outQueue_3_io_enq_bits),
    .io_deq_ready(outQueue_3_io_deq_ready),
    .io_deq_valid(outQueue_3_io_deq_valid),
    .io_deq_bits(outQueue_3_io_deq_bits)
  );
  Queue outQueue_4 ( // @[CGRAFullMask.scala 16:52]
    .clock(outQueue_4_clock),
    .reset(outQueue_4_reset),
    .io_enq_ready(outQueue_4_io_enq_ready),
    .io_enq_valid(outQueue_4_io_enq_valid),
    .io_enq_bits(outQueue_4_io_enq_bits),
    .io_deq_ready(outQueue_4_io_deq_ready),
    .io_deq_valid(outQueue_4_io_deq_valid),
    .io_deq_bits(outQueue_4_io_deq_bits)
  );
  Queue outQueue_5 ( // @[CGRAFullMask.scala 16:52]
    .clock(outQueue_5_clock),
    .reset(outQueue_5_reset),
    .io_enq_ready(outQueue_5_io_enq_ready),
    .io_enq_valid(outQueue_5_io_enq_valid),
    .io_enq_bits(outQueue_5_io_enq_bits),
    .io_deq_ready(outQueue_5_io_deq_ready),
    .io_deq_valid(outQueue_5_io_deq_valid),
    .io_deq_bits(outQueue_5_io_deq_bits)
  );
  Queue outQueue_6 ( // @[CGRAFullMask.scala 16:52]
    .clock(outQueue_6_clock),
    .reset(outQueue_6_reset),
    .io_enq_ready(outQueue_6_io_enq_ready),
    .io_enq_valid(outQueue_6_io_enq_valid),
    .io_enq_bits(outQueue_6_io_enq_bits),
    .io_deq_ready(outQueue_6_io_deq_ready),
    .io_deq_valid(outQueue_6_io_deq_valid),
    .io_deq_bits(outQueue_6_io_deq_bits)
  );
  Queue outQueue_7 ( // @[CGRAFullMask.scala 16:52]
    .clock(outQueue_7_clock),
    .reset(outQueue_7_reset),
    .io_enq_ready(outQueue_7_io_enq_ready),
    .io_enq_valid(outQueue_7_io_enq_valid),
    .io_enq_bits(outQueue_7_io_enq_bits),
    .io_deq_ready(outQueue_7_io_deq_ready),
    .io_deq_valid(outQueue_7_io_deq_valid),
    .io_deq_bits(outQueue_7_io_deq_bits)
  );
  Queue outQueue_8 ( // @[CGRAFullMask.scala 16:52]
    .clock(outQueue_8_clock),
    .reset(outQueue_8_reset),
    .io_enq_ready(outQueue_8_io_enq_ready),
    .io_enq_valid(outQueue_8_io_enq_valid),
    .io_enq_bits(outQueue_8_io_enq_bits),
    .io_deq_ready(outQueue_8_io_deq_ready),
    .io_deq_valid(outQueue_8_io_deq_valid),
    .io_deq_bits(outQueue_8_io_deq_bits)
  );
  Queue outQueue_9 ( // @[CGRAFullMask.scala 16:52]
    .clock(outQueue_9_clock),
    .reset(outQueue_9_reset),
    .io_enq_ready(outQueue_9_io_enq_ready),
    .io_enq_valid(outQueue_9_io_enq_valid),
    .io_enq_bits(outQueue_9_io_enq_bits),
    .io_deq_ready(outQueue_9_io_deq_ready),
    .io_deq_valid(outQueue_9_io_deq_valid),
    .io_deq_bits(outQueue_9_io_deq_bits)
  );
  Queue outQueue_10 ( // @[CGRAFullMask.scala 16:52]
    .clock(outQueue_10_clock),
    .reset(outQueue_10_reset),
    .io_enq_ready(outQueue_10_io_enq_ready),
    .io_enq_valid(outQueue_10_io_enq_valid),
    .io_enq_bits(outQueue_10_io_enq_bits),
    .io_deq_ready(outQueue_10_io_deq_ready),
    .io_deq_valid(outQueue_10_io_deq_valid),
    .io_deq_bits(outQueue_10_io_deq_bits)
  );
  Queue outQueue_11 ( // @[CGRAFullMask.scala 16:52]
    .clock(outQueue_11_clock),
    .reset(outQueue_11_reset),
    .io_enq_ready(outQueue_11_io_enq_ready),
    .io_enq_valid(outQueue_11_io_enq_valid),
    .io_enq_bits(outQueue_11_io_enq_bits),
    .io_deq_ready(outQueue_11_io_deq_ready),
    .io_deq_valid(outQueue_11_io_deq_valid),
    .io_deq_bits(outQueue_11_io_deq_bits)
  );
  Queue outQueue_12 ( // @[CGRAFullMask.scala 16:52]
    .clock(outQueue_12_clock),
    .reset(outQueue_12_reset),
    .io_enq_ready(outQueue_12_io_enq_ready),
    .io_enq_valid(outQueue_12_io_enq_valid),
    .io_enq_bits(outQueue_12_io_enq_bits),
    .io_deq_ready(outQueue_12_io_deq_ready),
    .io_deq_valid(outQueue_12_io_deq_valid),
    .io_deq_bits(outQueue_12_io_deq_bits)
  );
  Queue outQueue_13 ( // @[CGRAFullMask.scala 16:52]
    .clock(outQueue_13_clock),
    .reset(outQueue_13_reset),
    .io_enq_ready(outQueue_13_io_enq_ready),
    .io_enq_valid(outQueue_13_io_enq_valid),
    .io_enq_bits(outQueue_13_io_enq_bits),
    .io_deq_ready(outQueue_13_io_deq_ready),
    .io_deq_valid(outQueue_13_io_deq_valid),
    .io_deq_bits(outQueue_13_io_deq_bits)
  );
  Queue outQueue_14 ( // @[CGRAFullMask.scala 16:52]
    .clock(outQueue_14_clock),
    .reset(outQueue_14_reset),
    .io_enq_ready(outQueue_14_io_enq_ready),
    .io_enq_valid(outQueue_14_io_enq_valid),
    .io_enq_bits(outQueue_14_io_enq_bits),
    .io_deq_ready(outQueue_14_io_deq_ready),
    .io_deq_valid(outQueue_14_io_deq_valid),
    .io_deq_bits(outQueue_14_io_deq_bits)
  );
  Queue outQueue_15 ( // @[CGRAFullMask.scala 16:52]
    .clock(outQueue_15_clock),
    .reset(outQueue_15_reset),
    .io_enq_ready(outQueue_15_io_enq_ready),
    .io_enq_valid(outQueue_15_io_enq_valid),
    .io_enq_bits(outQueue_15_io_enq_bits),
    .io_deq_ready(outQueue_15_io_deq_ready),
    .io_deq_valid(outQueue_15_io_deq_valid),
    .io_deq_bits(outQueue_15_io_deq_bits)
  );
  SynInMask synInInst ( // @[CGRAFullMask.scala 19:25]
    .clock(synInInst_clock),
    .reset(synInInst_reset),
    .io_valid(synInInst_io_valid),
    .io_ready(synInInst_io_ready),
    .io_dataIn(synInInst_io_dataIn),
    .io_dataOut_0(synInInst_io_dataOut_0),
    .io_dataOut_1(synInInst_io_dataOut_1),
    .io_dataOut_2(synInInst_io_dataOut_2),
    .io_dataOut_3(synInInst_io_dataOut_3),
    .io_dataOut_4(synInInst_io_dataOut_4),
    .io_dataOut_5(synInInst_io_dataOut_5),
    .io_dataOut_6(synInInst_io_dataOut_6),
    .io_dataOut_7(synInInst_io_dataOut_7),
    .io_dataOut_8(synInInst_io_dataOut_8),
    .io_dataOut_9(synInInst_io_dataOut_9),
    .io_dataOut_10(synInInst_io_dataOut_10),
    .io_dataOut_11(synInInst_io_dataOut_11),
    .io_dataOut_12(synInInst_io_dataOut_12),
    .io_dataOut_13(synInInst_io_dataOut_13),
    .io_dataOut_14(synInInst_io_dataOut_14),
    .io_dataOut_15(synInInst_io_dataOut_15),
    .io_delayen(synInInst_io_delayen),
    .io_delayCycle(synInInst_io_delayCycle),
    .dmaEnWR_0(synInInst_dmaEnWR_0),
    .dmaCtrl_0(synInInst_dmaCtrl_0)
  );
  CGRAJ cgraInst ( // @[CGRAFullMask.scala 23:35]
    .clock(cgraInst_clock),
    .reset(cgraInst_reset),
    .io_cfgEn(cgraInst_io_cfgEn),
    .io_cfgAddr(cgraInst_io_cfgAddr),
    .io_cfgData(cgraInst_io_cfgData),
    .io_inputs_0(cgraInst_io_inputs_0),
    .io_inputs_1(cgraInst_io_inputs_1),
    .io_inputs_2(cgraInst_io_inputs_2),
    .io_inputs_3(cgraInst_io_inputs_3),
    .io_inputs_4(cgraInst_io_inputs_4),
    .io_inputs_5(cgraInst_io_inputs_5),
    .io_inputs_6(cgraInst_io_inputs_6),
    .io_inputs_7(cgraInst_io_inputs_7),
    .io_inputs_8(cgraInst_io_inputs_8),
    .io_inputs_9(cgraInst_io_inputs_9),
    .io_inputs_10(cgraInst_io_inputs_10),
    .io_inputs_11(cgraInst_io_inputs_11),
    .io_inputs_12(cgraInst_io_inputs_12),
    .io_inputs_13(cgraInst_io_inputs_13),
    .io_inputs_14(cgraInst_io_inputs_14),
    .io_inputs_15(cgraInst_io_inputs_15),
    .io_outputs_0(cgraInst_io_outputs_0),
    .io_outputs_1(cgraInst_io_outputs_1),
    .io_outputs_2(cgraInst_io_outputs_2),
    .io_outputs_3(cgraInst_io_outputs_3),
    .io_outputs_4(cgraInst_io_outputs_4),
    .io_outputs_5(cgraInst_io_outputs_5),
    .io_outputs_6(cgraInst_io_outputs_6),
    .io_outputs_7(cgraInst_io_outputs_7),
    .io_outputs_8(cgraInst_io_outputs_8),
    .io_outputs_9(cgraInst_io_outputs_9),
    .io_outputs_10(cgraInst_io_outputs_10),
    .io_outputs_11(cgraInst_io_outputs_11),
    .io_outputs_12(cgraInst_io_outputs_12),
    .io_outputs_13(cgraInst_io_outputs_13),
    .io_outputs_14(cgraInst_io_outputs_14),
    .io_outputs_15(cgraInst_io_outputs_15)
  );
  assign io_CGRAIO_ready = _T_143 | oneHot_18; // @[CGRAFullMask.scala 55:21]
  assign io_CGRAIO_data_read = {{32'd0}, _T_252}; // @[CGRAFullMask.scala 82:23]
  assign io_outputs_0 = cgraInst_io_outputs_0; // @[CGRAFullMask.scala 30:19]
  assign io_outputs_1 = cgraInst_io_outputs_1; // @[CGRAFullMask.scala 30:19]
  assign io_outputs_2 = cgraInst_io_outputs_2; // @[CGRAFullMask.scala 30:19]
  assign io_outputs_3 = cgraInst_io_outputs_3; // @[CGRAFullMask.scala 30:19]
  assign io_outputs_4 = cgraInst_io_outputs_4; // @[CGRAFullMask.scala 30:19]
  assign io_outputs_5 = cgraInst_io_outputs_5; // @[CGRAFullMask.scala 30:19]
  assign io_outputs_6 = cgraInst_io_outputs_6; // @[CGRAFullMask.scala 30:19]
  assign io_outputs_7 = cgraInst_io_outputs_7; // @[CGRAFullMask.scala 30:19]
  assign io_outputs_8 = cgraInst_io_outputs_8; // @[CGRAFullMask.scala 30:19]
  assign io_outputs_9 = cgraInst_io_outputs_9; // @[CGRAFullMask.scala 30:19]
  assign io_outputs_10 = cgraInst_io_outputs_10; // @[CGRAFullMask.scala 30:19]
  assign io_outputs_11 = cgraInst_io_outputs_11; // @[CGRAFullMask.scala 30:19]
  assign io_outputs_12 = cgraInst_io_outputs_12; // @[CGRAFullMask.scala 30:19]
  assign io_outputs_13 = cgraInst_io_outputs_13; // @[CGRAFullMask.scala 30:19]
  assign io_outputs_14 = cgraInst_io_outputs_14; // @[CGRAFullMask.scala 30:19]
  assign io_outputs_15 = cgraInst_io_outputs_15; // @[CGRAFullMask.scala 30:19]
  assign outQueue_0_clock = clock;
  assign outQueue_0_reset = reset;
  assign outQueue_0_io_enq_valid = cgraInst_io_outputs_0[32]; // @[CGRAFullMask.scala 29:30]
  assign outQueue_0_io_enq_bits = cgraInst_io_outputs_0[31:0]; // @[CGRAFullMask.scala 28:29]
  assign outQueue_0_io_deq_ready = _T_150 & io_CGRAIO_valid; // @[CGRAFullMask.scala 67:35]
  assign outQueue_1_clock = clock;
  assign outQueue_1_reset = reset;
  assign outQueue_1_io_enq_valid = cgraInst_io_outputs_1[32]; // @[CGRAFullMask.scala 29:30]
  assign outQueue_1_io_enq_bits = cgraInst_io_outputs_1[31:0]; // @[CGRAFullMask.scala 28:29]
  assign outQueue_1_io_deq_ready = _T_154 & io_CGRAIO_valid; // @[CGRAFullMask.scala 67:35]
  assign outQueue_2_clock = clock;
  assign outQueue_2_reset = reset;
  assign outQueue_2_io_enq_valid = cgraInst_io_outputs_2[32]; // @[CGRAFullMask.scala 29:30]
  assign outQueue_2_io_enq_bits = cgraInst_io_outputs_2[31:0]; // @[CGRAFullMask.scala 28:29]
  assign outQueue_2_io_deq_ready = _T_158 & io_CGRAIO_valid; // @[CGRAFullMask.scala 67:35]
  assign outQueue_3_clock = clock;
  assign outQueue_3_reset = reset;
  assign outQueue_3_io_enq_valid = cgraInst_io_outputs_3[32]; // @[CGRAFullMask.scala 29:30]
  assign outQueue_3_io_enq_bits = cgraInst_io_outputs_3[31:0]; // @[CGRAFullMask.scala 28:29]
  assign outQueue_3_io_deq_ready = _T_162 & io_CGRAIO_valid; // @[CGRAFullMask.scala 67:35]
  assign outQueue_4_clock = clock;
  assign outQueue_4_reset = reset;
  assign outQueue_4_io_enq_valid = cgraInst_io_outputs_4[32]; // @[CGRAFullMask.scala 29:30]
  assign outQueue_4_io_enq_bits = cgraInst_io_outputs_4[31:0]; // @[CGRAFullMask.scala 28:29]
  assign outQueue_4_io_deq_ready = _T_166 & io_CGRAIO_valid; // @[CGRAFullMask.scala 67:35]
  assign outQueue_5_clock = clock;
  assign outQueue_5_reset = reset;
  assign outQueue_5_io_enq_valid = cgraInst_io_outputs_5[32]; // @[CGRAFullMask.scala 29:30]
  assign outQueue_5_io_enq_bits = cgraInst_io_outputs_5[31:0]; // @[CGRAFullMask.scala 28:29]
  assign outQueue_5_io_deq_ready = _T_170 & io_CGRAIO_valid; // @[CGRAFullMask.scala 67:35]
  assign outQueue_6_clock = clock;
  assign outQueue_6_reset = reset;
  assign outQueue_6_io_enq_valid = cgraInst_io_outputs_6[32]; // @[CGRAFullMask.scala 29:30]
  assign outQueue_6_io_enq_bits = cgraInst_io_outputs_6[31:0]; // @[CGRAFullMask.scala 28:29]
  assign outQueue_6_io_deq_ready = _T_174 & io_CGRAIO_valid; // @[CGRAFullMask.scala 67:35]
  assign outQueue_7_clock = clock;
  assign outQueue_7_reset = reset;
  assign outQueue_7_io_enq_valid = cgraInst_io_outputs_7[32]; // @[CGRAFullMask.scala 29:30]
  assign outQueue_7_io_enq_bits = cgraInst_io_outputs_7[31:0]; // @[CGRAFullMask.scala 28:29]
  assign outQueue_7_io_deq_ready = _T_178 & io_CGRAIO_valid; // @[CGRAFullMask.scala 67:35]
  assign outQueue_8_clock = clock;
  assign outQueue_8_reset = reset;
  assign outQueue_8_io_enq_valid = cgraInst_io_outputs_8[32]; // @[CGRAFullMask.scala 29:30]
  assign outQueue_8_io_enq_bits = cgraInst_io_outputs_8[31:0]; // @[CGRAFullMask.scala 28:29]
  assign outQueue_8_io_deq_ready = _T_182 & io_CGRAIO_valid; // @[CGRAFullMask.scala 67:35]
  assign outQueue_9_clock = clock;
  assign outQueue_9_reset = reset;
  assign outQueue_9_io_enq_valid = cgraInst_io_outputs_9[32]; // @[CGRAFullMask.scala 29:30]
  assign outQueue_9_io_enq_bits = cgraInst_io_outputs_9[31:0]; // @[CGRAFullMask.scala 28:29]
  assign outQueue_9_io_deq_ready = _T_186 & io_CGRAIO_valid; // @[CGRAFullMask.scala 67:35]
  assign outQueue_10_clock = clock;
  assign outQueue_10_reset = reset;
  assign outQueue_10_io_enq_valid = cgraInst_io_outputs_10[32]; // @[CGRAFullMask.scala 29:30]
  assign outQueue_10_io_enq_bits = cgraInst_io_outputs_10[31:0]; // @[CGRAFullMask.scala 28:29]
  assign outQueue_10_io_deq_ready = _T_190 & io_CGRAIO_valid; // @[CGRAFullMask.scala 67:35]
  assign outQueue_11_clock = clock;
  assign outQueue_11_reset = reset;
  assign outQueue_11_io_enq_valid = cgraInst_io_outputs_11[32]; // @[CGRAFullMask.scala 29:30]
  assign outQueue_11_io_enq_bits = cgraInst_io_outputs_11[31:0]; // @[CGRAFullMask.scala 28:29]
  assign outQueue_11_io_deq_ready = _T_194 & io_CGRAIO_valid; // @[CGRAFullMask.scala 67:35]
  assign outQueue_12_clock = clock;
  assign outQueue_12_reset = reset;
  assign outQueue_12_io_enq_valid = cgraInst_io_outputs_12[32]; // @[CGRAFullMask.scala 29:30]
  assign outQueue_12_io_enq_bits = cgraInst_io_outputs_12[31:0]; // @[CGRAFullMask.scala 28:29]
  assign outQueue_12_io_deq_ready = _T_198 & io_CGRAIO_valid; // @[CGRAFullMask.scala 67:35]
  assign outQueue_13_clock = clock;
  assign outQueue_13_reset = reset;
  assign outQueue_13_io_enq_valid = cgraInst_io_outputs_13[32]; // @[CGRAFullMask.scala 29:30]
  assign outQueue_13_io_enq_bits = cgraInst_io_outputs_13[31:0]; // @[CGRAFullMask.scala 28:29]
  assign outQueue_13_io_deq_ready = _T_202 & io_CGRAIO_valid; // @[CGRAFullMask.scala 67:35]
  assign outQueue_14_clock = clock;
  assign outQueue_14_reset = reset;
  assign outQueue_14_io_enq_valid = cgraInst_io_outputs_14[32]; // @[CGRAFullMask.scala 29:30]
  assign outQueue_14_io_enq_bits = cgraInst_io_outputs_14[31:0]; // @[CGRAFullMask.scala 28:29]
  assign outQueue_14_io_deq_ready = _T_206 & io_CGRAIO_valid; // @[CGRAFullMask.scala 67:35]
  assign outQueue_15_clock = clock;
  assign outQueue_15_reset = reset;
  assign outQueue_15_io_enq_valid = cgraInst_io_outputs_15[32]; // @[CGRAFullMask.scala 29:30]
  assign outQueue_15_io_enq_bits = cgraInst_io_outputs_15[31:0]; // @[CGRAFullMask.scala 28:29]
  assign outQueue_15_io_deq_ready = _T_210 & io_CGRAIO_valid; // @[CGRAFullMask.scala 67:35]
  assign synInInst_clock = clock;
  assign synInInst_reset = reset;
  assign synInInst_io_valid = _T_146 & addrIsW; // @[CGRAFullMask.scala 65:22]
  assign synInInst_io_dataIn = io_CGRAIO_data_write; // @[CGRAFullMask.scala 77:23]
  assign synInInst_io_delayen = _T_218 & io_CGRAIO_valid; // @[CGRAFullMask.scala 70:24]
  assign synInInst_io_delayCycle = io_CGRAIO_data_write; // @[CGRAFullMask.scala 80:27]
  assign synInInst_dmaEnWR_0 = _T_100_0;
  assign synInInst_dmaCtrl_0 = dmaCtrl;
  assign cgraInst_clock = clock;
  assign cgraInst_reset = reset;
  assign cgraInst_io_cfgEn = _T_214 & io_CGRAIO_valid; // @[CGRAFullMask.scala 69:21]
  assign cgraInst_io_cfgAddr = io_CGRAIO_data_write[40:32]; // @[CGRAFullMask.scala 79:23]
  assign cgraInst_io_cfgData = io_CGRAIO_data_write[31:0]; // @[CGRAFullMask.scala 78:23]
  assign cgraInst_io_inputs_0 = synInInst_io_dataOut_0; // @[CGRAFullMask.scala 27:27]
  assign cgraInst_io_inputs_1 = synInInst_io_dataOut_1; // @[CGRAFullMask.scala 27:27]
  assign cgraInst_io_inputs_2 = synInInst_io_dataOut_2; // @[CGRAFullMask.scala 27:27]
  assign cgraInst_io_inputs_3 = synInInst_io_dataOut_3; // @[CGRAFullMask.scala 27:27]
  assign cgraInst_io_inputs_4 = synInInst_io_dataOut_4; // @[CGRAFullMask.scala 27:27]
  assign cgraInst_io_inputs_5 = synInInst_io_dataOut_5; // @[CGRAFullMask.scala 27:27]
  assign cgraInst_io_inputs_6 = synInInst_io_dataOut_6; // @[CGRAFullMask.scala 27:27]
  assign cgraInst_io_inputs_7 = synInInst_io_dataOut_7; // @[CGRAFullMask.scala 27:27]
  assign cgraInst_io_inputs_8 = synInInst_io_dataOut_8; // @[CGRAFullMask.scala 27:27]
  assign cgraInst_io_inputs_9 = synInInst_io_dataOut_9; // @[CGRAFullMask.scala 27:27]
  assign cgraInst_io_inputs_10 = synInInst_io_dataOut_10; // @[CGRAFullMask.scala 27:27]
  assign cgraInst_io_inputs_11 = synInInst_io_dataOut_11; // @[CGRAFullMask.scala 27:27]
  assign cgraInst_io_inputs_12 = synInInst_io_dataOut_12; // @[CGRAFullMask.scala 27:27]
  assign cgraInst_io_inputs_13 = synInInst_io_dataOut_13; // @[CGRAFullMask.scala 27:27]
  assign cgraInst_io_inputs_14 = synInInst_io_dataOut_14; // @[CGRAFullMask.scala 27:27]
  assign cgraInst_io_inputs_15 = synInInst_io_dataOut_15; // @[CGRAFullMask.scala 27:27]
endmodule
module iFetch(
  input         clock,
  input         reset,
  input  [31:0] io_instIn,
  output [31:0] io_instOut,
  output [31:0] io_pc,
  output [31:0] io_snpc,
  input  [31:0] io_dnpc,
  input         io_jump,
  input         intrTimeCnt_0,
  input         hazardPCBlock_0,
  input         blockDMA_0,
  input         block23_0,
  input         block1_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] pc; // @[Reg.scala 27:20]
  wire [31:0] snpc = pc + 32'h4; // @[iFetch.scala 41:14]
  wire  _T_1 = block1_0 | block23_0; // @[iFetch.scala 39:78]
  wire  _T_2 = _T_1 | blockDMA_0; // @[iFetch.scala 39:88]
  wire  _T_3 = ~_T_2; // @[iFetch.scala 39:70]
  wire  _T_4 = ~hazardPCBlock_0; // @[iFetch.scala 39:105]
  wire  _T_5 = _T_4 | intrTimeCnt_0; // @[iFetch.scala 39:120]
  wire  _T_6 = _T_3 & _T_5; // @[iFetch.scala 39:101]
  assign io_instOut = io_instIn; // @[iFetch.scala 56:14]
  assign io_pc = pc; // @[iFetch.scala 49:9]
  assign io_snpc = pc + 32'h4; // @[iFetch.scala 42:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pc <= 32'h80000000;
    end else if (_T_6) begin
      if (io_jump) begin
        pc <= io_dnpc;
      end else begin
        pc <= snpc;
      end
    end
  end
endmodule
module immeGen(
  input  [31:0] io_inst,
  output [63:0] io_imme
);
  wire [51:0] _T_3 = io_inst[31] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] Iimm = {_T_3,io_inst[31:20]}; // @[Cat.scala 29:58]
  wire [11:0] _T_6 = {io_inst[31:25],io_inst[11:7]}; // @[Cat.scala 29:58]
  wire [51:0] _T_9 = _T_6[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] Simm = {_T_9,io_inst[31:25],io_inst[11:7]}; // @[Cat.scala 29:58]
  wire [12:0] _T_17 = {io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8],1'h0}; // @[Cat.scala 29:58]
  wire [50:0] _T_20 = _T_17[12] ? 51'h7ffffffffffff : 51'h0; // @[Bitwise.scala 72:12]
  wire [63:0] Bimm = {_T_20,io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_22 = {io_inst[31:12],12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_25 = _T_22[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] Uimm = {_T_25,io_inst[31:12],12'h0}; // @[Cat.scala 29:58]
  wire [20:0] _T_33 = {io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21],1'h0}; // @[Cat.scala 29:58]
  wire [42:0] _T_36 = _T_33[20] ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 72:12]
  wire [63:0] Jimm = {_T_36,io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_37 = io_inst & 32'h707f; // @[immeGen.scala 55:47]
  wire  _T_38 = 32'h3023 == _T_37; // @[immeGen.scala 55:47]
  wire [31:0] _T_39 = io_inst & 32'hfc00707f; // @[immeGen.scala 52:47]
  wire  _T_40 = 32'h1013 == _T_39; // @[immeGen.scala 52:47]
  wire  _T_42 = 32'h6063 == _T_37; // @[immeGen.scala 56:47]
  wire  _T_44 = 32'h1003 == _T_37; // @[immeGen.scala 52:47]
  wire  _T_46 = 32'h4013 == _T_37; // @[immeGen.scala 52:47]
  wire [31:0] _T_47 = io_inst & 32'h7f; // @[immeGen.scala 53:47]
  wire  _T_48 = 32'h6f == _T_47; // @[immeGen.scala 53:47]
  wire  _T_50 = 32'h6013 == _T_37; // @[immeGen.scala 52:47]
  wire  _T_52 = 32'h5063 == _T_37; // @[immeGen.scala 56:47]
  wire  _T_54 = 32'h7013 == _T_37; // @[immeGen.scala 52:47]
  wire  _T_56 = 32'h4003 == _T_37; // @[immeGen.scala 52:47]
  wire  _T_58 = 32'h3 == _T_37; // @[immeGen.scala 52:47]
  wire  _T_60 = 32'h2023 == _T_37; // @[immeGen.scala 55:47]
  wire  _T_62 = 32'h1063 == _T_37; // @[immeGen.scala 56:47]
  wire  _T_64 = 32'h1b == _T_37; // @[immeGen.scala 52:47]
  wire  _T_66 = 32'h17 == _T_47; // @[immeGen.scala 54:47]
  wire  _T_68 = 32'h4063 == _T_37; // @[immeGen.scala 56:47]
  wire  _T_70 = 32'h40005013 == _T_39; // @[immeGen.scala 52:47]
  wire  _T_72 = 32'h63 == _T_37; // @[immeGen.scala 56:47]
  wire  _T_74 = 32'h3003 == _T_37; // @[immeGen.scala 52:47]
  wire [31:0] _T_75 = io_inst & 32'hfe00707f; // @[immeGen.scala 52:47]
  wire  _T_76 = 32'h4000501b == _T_75; // @[immeGen.scala 52:47]
  wire  _T_78 = 32'h67 == _T_37; // @[immeGen.scala 52:47]
  wire  _T_80 = 32'h5013 == _T_39; // @[immeGen.scala 52:47]
  wire  _T_82 = 32'h23 == _T_37; // @[immeGen.scala 55:47]
  wire  _T_84 = 32'h37 == _T_47; // @[immeGen.scala 54:47]
  wire  _T_86 = 32'h501b == _T_75; // @[immeGen.scala 52:47]
  wire  _T_88 = 32'h5003 == _T_37; // @[immeGen.scala 52:47]
  wire  _T_90 = 32'h6003 == _T_37; // @[immeGen.scala 52:47]
  wire  _T_92 = 32'h2003 == _T_37; // @[immeGen.scala 52:47]
  wire  _T_94 = 32'h101b == _T_75; // @[immeGen.scala 52:47]
  wire  _T_96 = 32'h1023 == _T_37; // @[immeGen.scala 55:47]
  wire  _T_98 = 32'h13 == _T_37; // @[immeGen.scala 52:47]
  wire  _T_100 = 32'h7063 == _T_37; // @[immeGen.scala 56:47]
  wire  _T_102 = 32'h3013 == _T_37; // @[immeGen.scala 52:47]
  wire  _T_104 = 32'h1073 == _T_37; // @[immeGen.scala 62:29]
  wire  _T_106 = 32'h2073 == _T_37; // @[immeGen.scala 63:29]
  wire  _T_108 = 32'h6073 == _T_37; // @[immeGen.scala 64:29]
  wire  _T_110 = 32'h7073 == _T_37; // @[immeGen.scala 65:29]
  wire  _T_112 = 32'h3073 == _T_37; // @[immeGen.scala 66:29]
  wire [63:0] _T_113 = _T_112 ? Iimm : 64'h0; // @[Mux.scala 98:16]
  wire [63:0] _T_114 = _T_110 ? Iimm : _T_113; // @[Mux.scala 98:16]
  wire [63:0] _T_115 = _T_108 ? Iimm : _T_114; // @[Mux.scala 98:16]
  wire [63:0] _T_116 = _T_106 ? Iimm : _T_115; // @[Mux.scala 98:16]
  wire [63:0] _T_117 = _T_104 ? Iimm : _T_116; // @[Mux.scala 98:16]
  wire [63:0] _T_118 = _T_102 ? Iimm : _T_117; // @[Mux.scala 98:16]
  wire [63:0] _T_119 = _T_100 ? Bimm : _T_118; // @[Mux.scala 98:16]
  wire [63:0] _T_120 = _T_98 ? Iimm : _T_119; // @[Mux.scala 98:16]
  wire [63:0] _T_121 = _T_96 ? Simm : _T_120; // @[Mux.scala 98:16]
  wire [63:0] _T_122 = _T_94 ? Iimm : _T_121; // @[Mux.scala 98:16]
  wire [63:0] _T_123 = _T_92 ? Iimm : _T_122; // @[Mux.scala 98:16]
  wire [63:0] _T_124 = _T_90 ? Iimm : _T_123; // @[Mux.scala 98:16]
  wire [63:0] _T_125 = _T_88 ? Iimm : _T_124; // @[Mux.scala 98:16]
  wire [63:0] _T_126 = _T_86 ? Iimm : _T_125; // @[Mux.scala 98:16]
  wire [63:0] _T_127 = _T_84 ? Uimm : _T_126; // @[Mux.scala 98:16]
  wire [63:0] _T_128 = _T_82 ? Simm : _T_127; // @[Mux.scala 98:16]
  wire [63:0] _T_129 = _T_80 ? Iimm : _T_128; // @[Mux.scala 98:16]
  wire [63:0] _T_130 = _T_78 ? Iimm : _T_129; // @[Mux.scala 98:16]
  wire [63:0] _T_131 = _T_76 ? Iimm : _T_130; // @[Mux.scala 98:16]
  wire [63:0] _T_132 = _T_74 ? Iimm : _T_131; // @[Mux.scala 98:16]
  wire [63:0] _T_133 = _T_72 ? Bimm : _T_132; // @[Mux.scala 98:16]
  wire [63:0] _T_134 = _T_70 ? Iimm : _T_133; // @[Mux.scala 98:16]
  wire [63:0] _T_135 = _T_68 ? Bimm : _T_134; // @[Mux.scala 98:16]
  wire [63:0] _T_136 = _T_66 ? Uimm : _T_135; // @[Mux.scala 98:16]
  wire [63:0] _T_137 = _T_64 ? Iimm : _T_136; // @[Mux.scala 98:16]
  wire [63:0] _T_138 = _T_62 ? Bimm : _T_137; // @[Mux.scala 98:16]
  wire [63:0] _T_139 = _T_60 ? Simm : _T_138; // @[Mux.scala 98:16]
  wire [63:0] _T_140 = _T_58 ? Iimm : _T_139; // @[Mux.scala 98:16]
  wire [63:0] _T_141 = _T_56 ? Iimm : _T_140; // @[Mux.scala 98:16]
  wire [63:0] _T_142 = _T_54 ? Iimm : _T_141; // @[Mux.scala 98:16]
  wire [63:0] _T_143 = _T_52 ? Bimm : _T_142; // @[Mux.scala 98:16]
  wire [63:0] _T_144 = _T_50 ? Iimm : _T_143; // @[Mux.scala 98:16]
  wire [63:0] _T_145 = _T_48 ? Jimm : _T_144; // @[Mux.scala 98:16]
  wire [63:0] _T_146 = _T_46 ? Iimm : _T_145; // @[Mux.scala 98:16]
  wire [63:0] _T_147 = _T_44 ? Iimm : _T_146; // @[Mux.scala 98:16]
  wire [63:0] _T_148 = _T_42 ? Bimm : _T_147; // @[Mux.scala 98:16]
  wire [63:0] _T_149 = _T_40 ? Iimm : _T_148; // @[Mux.scala 98:16]
  assign io_imme = _T_38 ? Simm : _T_149; // @[immeGen.scala 68:13]
endmodule
module RF(
  input         clock,
  input         reset,
  input  [31:0] io_pc,
  input         io_we,
  input  [4:0]  io_rs1,
  input  [4:0]  io_rs2,
  input  [4:0]  io_rd,
  input  [4:0]  io_rdID,
  output [63:0] io_dout1,
  output [63:0] io_dout2,
  output [63:0] io_rdDout,
  input  [63:0] io_din,
  output [63:0] io_doutWB,
  input         blockDMA_0,
  input         block23_0,
  input         block1_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] DPIC_RegRead_ins_inst_0; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_1; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_2; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_3; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_4; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_5; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_6; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_7; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_8; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_9; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_10; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_11; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_12; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_13; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_14; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_15; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_16; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_17; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_18; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_19; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_20; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_21; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_22; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_23; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_24; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_25; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_26; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_27; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_28; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_29; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_30; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_inst_31; // @[regFile.scala 30:33]
  wire [63:0] DPIC_RegRead_ins_pc; // @[regFile.scala 30:33]
  wire  _T_1 = block1_0 | block23_0; // @[regFile.scala 57:50]
  wire  _T_2 = _T_1 | blockDMA_0; // @[regFile.scala 57:61]
  wire  _T_3 = ~_T_2; // @[regFile.scala 57:41]
  wire  _T_7 = io_rd == 5'h1; // @[regFile.scala 55:22]
  wire  _T_8 = io_we & _T_7; // @[regFile.scala 55:13]
  wire  _T_12 = _T_8 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_13; // @[Reg.scala 15:16]
  wire  _T_15 = io_rd == 5'h2; // @[regFile.scala 55:22]
  wire  _T_16 = io_we & _T_15; // @[regFile.scala 55:13]
  wire  _T_20 = _T_16 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_21; // @[Reg.scala 15:16]
  wire  _T_23 = io_rd == 5'h3; // @[regFile.scala 55:22]
  wire  _T_24 = io_we & _T_23; // @[regFile.scala 55:13]
  wire  _T_28 = _T_24 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_29; // @[Reg.scala 15:16]
  wire  _T_31 = io_rd == 5'h4; // @[regFile.scala 55:22]
  wire  _T_32 = io_we & _T_31; // @[regFile.scala 55:13]
  wire  _T_36 = _T_32 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_37; // @[Reg.scala 15:16]
  wire  _T_39 = io_rd == 5'h5; // @[regFile.scala 55:22]
  wire  _T_40 = io_we & _T_39; // @[regFile.scala 55:13]
  wire  _T_44 = _T_40 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_45; // @[Reg.scala 15:16]
  wire  _T_47 = io_rd == 5'h6; // @[regFile.scala 55:22]
  wire  _T_48 = io_we & _T_47; // @[regFile.scala 55:13]
  wire  _T_52 = _T_48 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_53; // @[Reg.scala 15:16]
  wire  _T_55 = io_rd == 5'h7; // @[regFile.scala 55:22]
  wire  _T_56 = io_we & _T_55; // @[regFile.scala 55:13]
  wire  _T_60 = _T_56 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_61; // @[Reg.scala 15:16]
  wire  _T_63 = io_rd == 5'h8; // @[regFile.scala 55:22]
  wire  _T_64 = io_we & _T_63; // @[regFile.scala 55:13]
  wire  _T_68 = _T_64 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_69; // @[Reg.scala 15:16]
  wire  _T_71 = io_rd == 5'h9; // @[regFile.scala 55:22]
  wire  _T_72 = io_we & _T_71; // @[regFile.scala 55:13]
  wire  _T_76 = _T_72 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_77; // @[Reg.scala 15:16]
  wire  _T_79 = io_rd == 5'ha; // @[regFile.scala 55:22]
  wire  _T_80 = io_we & _T_79; // @[regFile.scala 55:13]
  wire  _T_84 = _T_80 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_85; // @[Reg.scala 15:16]
  wire  _T_87 = io_rd == 5'hb; // @[regFile.scala 55:22]
  wire  _T_88 = io_we & _T_87; // @[regFile.scala 55:13]
  wire  _T_92 = _T_88 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_93; // @[Reg.scala 15:16]
  wire  _T_95 = io_rd == 5'hc; // @[regFile.scala 55:22]
  wire  _T_96 = io_we & _T_95; // @[regFile.scala 55:13]
  wire  _T_100 = _T_96 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_101; // @[Reg.scala 15:16]
  wire  _T_103 = io_rd == 5'hd; // @[regFile.scala 55:22]
  wire  _T_104 = io_we & _T_103; // @[regFile.scala 55:13]
  wire  _T_108 = _T_104 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_109; // @[Reg.scala 15:16]
  wire  _T_111 = io_rd == 5'he; // @[regFile.scala 55:22]
  wire  _T_112 = io_we & _T_111; // @[regFile.scala 55:13]
  wire  _T_116 = _T_112 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_117; // @[Reg.scala 15:16]
  wire  _T_119 = io_rd == 5'hf; // @[regFile.scala 55:22]
  wire  _T_120 = io_we & _T_119; // @[regFile.scala 55:13]
  wire  _T_124 = _T_120 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_125; // @[Reg.scala 15:16]
  wire  _T_127 = io_rd == 5'h10; // @[regFile.scala 55:22]
  wire  _T_128 = io_we & _T_127; // @[regFile.scala 55:13]
  wire  _T_132 = _T_128 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_133; // @[Reg.scala 15:16]
  wire  _T_135 = io_rd == 5'h11; // @[regFile.scala 55:22]
  wire  _T_136 = io_we & _T_135; // @[regFile.scala 55:13]
  wire  _T_140 = _T_136 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_141; // @[Reg.scala 15:16]
  wire  _T_143 = io_rd == 5'h12; // @[regFile.scala 55:22]
  wire  _T_144 = io_we & _T_143; // @[regFile.scala 55:13]
  wire  _T_148 = _T_144 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_149; // @[Reg.scala 15:16]
  wire  _T_151 = io_rd == 5'h13; // @[regFile.scala 55:22]
  wire  _T_152 = io_we & _T_151; // @[regFile.scala 55:13]
  wire  _T_156 = _T_152 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_157; // @[Reg.scala 15:16]
  wire  _T_159 = io_rd == 5'h14; // @[regFile.scala 55:22]
  wire  _T_160 = io_we & _T_159; // @[regFile.scala 55:13]
  wire  _T_164 = _T_160 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_165; // @[Reg.scala 15:16]
  wire  _T_167 = io_rd == 5'h15; // @[regFile.scala 55:22]
  wire  _T_168 = io_we & _T_167; // @[regFile.scala 55:13]
  wire  _T_172 = _T_168 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_173; // @[Reg.scala 15:16]
  wire  _T_175 = io_rd == 5'h16; // @[regFile.scala 55:22]
  wire  _T_176 = io_we & _T_175; // @[regFile.scala 55:13]
  wire  _T_180 = _T_176 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_181; // @[Reg.scala 15:16]
  wire  _T_183 = io_rd == 5'h17; // @[regFile.scala 55:22]
  wire  _T_184 = io_we & _T_183; // @[regFile.scala 55:13]
  wire  _T_188 = _T_184 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_189; // @[Reg.scala 15:16]
  wire  _T_191 = io_rd == 5'h18; // @[regFile.scala 55:22]
  wire  _T_192 = io_we & _T_191; // @[regFile.scala 55:13]
  wire  _T_196 = _T_192 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_197; // @[Reg.scala 15:16]
  wire  _T_199 = io_rd == 5'h19; // @[regFile.scala 55:22]
  wire  _T_200 = io_we & _T_199; // @[regFile.scala 55:13]
  wire  _T_204 = _T_200 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_205; // @[Reg.scala 15:16]
  wire  _T_207 = io_rd == 5'h1a; // @[regFile.scala 55:22]
  wire  _T_208 = io_we & _T_207; // @[regFile.scala 55:13]
  wire  _T_212 = _T_208 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_213; // @[Reg.scala 15:16]
  wire  _T_215 = io_rd == 5'h1b; // @[regFile.scala 55:22]
  wire  _T_216 = io_we & _T_215; // @[regFile.scala 55:13]
  wire  _T_220 = _T_216 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_221; // @[Reg.scala 15:16]
  wire  _T_223 = io_rd == 5'h1c; // @[regFile.scala 55:22]
  wire  _T_224 = io_we & _T_223; // @[regFile.scala 55:13]
  wire  _T_228 = _T_224 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_229; // @[Reg.scala 15:16]
  wire  _T_231 = io_rd == 5'h1d; // @[regFile.scala 55:22]
  wire  _T_232 = io_we & _T_231; // @[regFile.scala 55:13]
  wire  _T_236 = _T_232 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_237; // @[Reg.scala 15:16]
  wire  _T_239 = io_rd == 5'h1e; // @[regFile.scala 55:22]
  wire  _T_240 = io_we & _T_239; // @[regFile.scala 55:13]
  wire  _T_244 = _T_240 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_245; // @[Reg.scala 15:16]
  wire  _T_247 = io_rd == 5'h1f; // @[regFile.scala 55:22]
  wire  _T_248 = io_we & _T_247; // @[regFile.scala 55:13]
  wire  _T_252 = _T_248 & _T_3; // @[regFile.scala 57:38]
  reg [63:0] _T_253; // @[Reg.scala 15:16]
  wire  _T_254 = 5'h1 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_255 = _T_254 ? _T_13 : 64'h0; // @[Mux.scala 80:57]
  wire  _T_256 = 5'h2 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_257 = _T_256 ? _T_21 : _T_255; // @[Mux.scala 80:57]
  wire  _T_258 = 5'h3 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_259 = _T_258 ? _T_29 : _T_257; // @[Mux.scala 80:57]
  wire  _T_260 = 5'h4 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_261 = _T_260 ? _T_37 : _T_259; // @[Mux.scala 80:57]
  wire  _T_262 = 5'h5 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_263 = _T_262 ? _T_45 : _T_261; // @[Mux.scala 80:57]
  wire  _T_264 = 5'h6 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_265 = _T_264 ? _T_53 : _T_263; // @[Mux.scala 80:57]
  wire  _T_266 = 5'h7 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_267 = _T_266 ? _T_61 : _T_265; // @[Mux.scala 80:57]
  wire  _T_268 = 5'h8 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_269 = _T_268 ? _T_69 : _T_267; // @[Mux.scala 80:57]
  wire  _T_270 = 5'h9 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_271 = _T_270 ? _T_77 : _T_269; // @[Mux.scala 80:57]
  wire  _T_272 = 5'ha == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_273 = _T_272 ? _T_85 : _T_271; // @[Mux.scala 80:57]
  wire  _T_274 = 5'hb == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_275 = _T_274 ? _T_93 : _T_273; // @[Mux.scala 80:57]
  wire  _T_276 = 5'hc == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_277 = _T_276 ? _T_101 : _T_275; // @[Mux.scala 80:57]
  wire  _T_278 = 5'hd == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_279 = _T_278 ? _T_109 : _T_277; // @[Mux.scala 80:57]
  wire  _T_280 = 5'he == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_281 = _T_280 ? _T_117 : _T_279; // @[Mux.scala 80:57]
  wire  _T_282 = 5'hf == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_283 = _T_282 ? _T_125 : _T_281; // @[Mux.scala 80:57]
  wire  _T_284 = 5'h10 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_285 = _T_284 ? _T_133 : _T_283; // @[Mux.scala 80:57]
  wire  _T_286 = 5'h11 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_287 = _T_286 ? _T_141 : _T_285; // @[Mux.scala 80:57]
  wire  _T_288 = 5'h12 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_289 = _T_288 ? _T_149 : _T_287; // @[Mux.scala 80:57]
  wire  _T_290 = 5'h13 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_291 = _T_290 ? _T_157 : _T_289; // @[Mux.scala 80:57]
  wire  _T_292 = 5'h14 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_293 = _T_292 ? _T_165 : _T_291; // @[Mux.scala 80:57]
  wire  _T_294 = 5'h15 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_295 = _T_294 ? _T_173 : _T_293; // @[Mux.scala 80:57]
  wire  _T_296 = 5'h16 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_297 = _T_296 ? _T_181 : _T_295; // @[Mux.scala 80:57]
  wire  _T_298 = 5'h17 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_299 = _T_298 ? _T_189 : _T_297; // @[Mux.scala 80:57]
  wire  _T_300 = 5'h18 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_301 = _T_300 ? _T_197 : _T_299; // @[Mux.scala 80:57]
  wire  _T_302 = 5'h19 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_303 = _T_302 ? _T_205 : _T_301; // @[Mux.scala 80:57]
  wire  _T_304 = 5'h1a == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_305 = _T_304 ? _T_213 : _T_303; // @[Mux.scala 80:57]
  wire  _T_306 = 5'h1b == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_307 = _T_306 ? _T_221 : _T_305; // @[Mux.scala 80:57]
  wire  _T_308 = 5'h1c == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_309 = _T_308 ? _T_229 : _T_307; // @[Mux.scala 80:57]
  wire  _T_310 = 5'h1d == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_311 = _T_310 ? _T_237 : _T_309; // @[Mux.scala 80:57]
  wire  _T_312 = 5'h1e == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_313 = _T_312 ? _T_245 : _T_311; // @[Mux.scala 80:57]
  wire  _T_314 = 5'h1f == io_rs1; // @[Mux.scala 80:60]
  wire  _T_316 = 5'h1 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_317 = _T_316 ? _T_13 : 64'h0; // @[Mux.scala 80:57]
  wire  _T_318 = 5'h2 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_319 = _T_318 ? _T_21 : _T_317; // @[Mux.scala 80:57]
  wire  _T_320 = 5'h3 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_321 = _T_320 ? _T_29 : _T_319; // @[Mux.scala 80:57]
  wire  _T_322 = 5'h4 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_323 = _T_322 ? _T_37 : _T_321; // @[Mux.scala 80:57]
  wire  _T_324 = 5'h5 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_325 = _T_324 ? _T_45 : _T_323; // @[Mux.scala 80:57]
  wire  _T_326 = 5'h6 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_327 = _T_326 ? _T_53 : _T_325; // @[Mux.scala 80:57]
  wire  _T_328 = 5'h7 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_329 = _T_328 ? _T_61 : _T_327; // @[Mux.scala 80:57]
  wire  _T_330 = 5'h8 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_331 = _T_330 ? _T_69 : _T_329; // @[Mux.scala 80:57]
  wire  _T_332 = 5'h9 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_333 = _T_332 ? _T_77 : _T_331; // @[Mux.scala 80:57]
  wire  _T_334 = 5'ha == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_335 = _T_334 ? _T_85 : _T_333; // @[Mux.scala 80:57]
  wire  _T_336 = 5'hb == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_337 = _T_336 ? _T_93 : _T_335; // @[Mux.scala 80:57]
  wire  _T_338 = 5'hc == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_339 = _T_338 ? _T_101 : _T_337; // @[Mux.scala 80:57]
  wire  _T_340 = 5'hd == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_341 = _T_340 ? _T_109 : _T_339; // @[Mux.scala 80:57]
  wire  _T_342 = 5'he == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_343 = _T_342 ? _T_117 : _T_341; // @[Mux.scala 80:57]
  wire  _T_344 = 5'hf == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_345 = _T_344 ? _T_125 : _T_343; // @[Mux.scala 80:57]
  wire  _T_346 = 5'h10 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_347 = _T_346 ? _T_133 : _T_345; // @[Mux.scala 80:57]
  wire  _T_348 = 5'h11 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_349 = _T_348 ? _T_141 : _T_347; // @[Mux.scala 80:57]
  wire  _T_350 = 5'h12 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_351 = _T_350 ? _T_149 : _T_349; // @[Mux.scala 80:57]
  wire  _T_352 = 5'h13 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_353 = _T_352 ? _T_157 : _T_351; // @[Mux.scala 80:57]
  wire  _T_354 = 5'h14 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_355 = _T_354 ? _T_165 : _T_353; // @[Mux.scala 80:57]
  wire  _T_356 = 5'h15 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_357 = _T_356 ? _T_173 : _T_355; // @[Mux.scala 80:57]
  wire  _T_358 = 5'h16 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_359 = _T_358 ? _T_181 : _T_357; // @[Mux.scala 80:57]
  wire  _T_360 = 5'h17 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_361 = _T_360 ? _T_189 : _T_359; // @[Mux.scala 80:57]
  wire  _T_362 = 5'h18 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_363 = _T_362 ? _T_197 : _T_361; // @[Mux.scala 80:57]
  wire  _T_364 = 5'h19 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_365 = _T_364 ? _T_205 : _T_363; // @[Mux.scala 80:57]
  wire  _T_366 = 5'h1a == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_367 = _T_366 ? _T_213 : _T_365; // @[Mux.scala 80:57]
  wire  _T_368 = 5'h1b == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_369 = _T_368 ? _T_221 : _T_367; // @[Mux.scala 80:57]
  wire  _T_370 = 5'h1c == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_371 = _T_370 ? _T_229 : _T_369; // @[Mux.scala 80:57]
  wire  _T_372 = 5'h1d == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_373 = _T_372 ? _T_237 : _T_371; // @[Mux.scala 80:57]
  wire  _T_374 = 5'h1e == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_375 = _T_374 ? _T_245 : _T_373; // @[Mux.scala 80:57]
  wire  _T_376 = 5'h1f == io_rs2; // @[Mux.scala 80:60]
  wire  _T_378 = 5'h1 == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_379 = _T_378 ? _T_13 : 64'h0; // @[Mux.scala 80:57]
  wire  _T_380 = 5'h2 == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_381 = _T_380 ? _T_21 : _T_379; // @[Mux.scala 80:57]
  wire  _T_382 = 5'h3 == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_383 = _T_382 ? _T_29 : _T_381; // @[Mux.scala 80:57]
  wire  _T_384 = 5'h4 == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_385 = _T_384 ? _T_37 : _T_383; // @[Mux.scala 80:57]
  wire  _T_386 = 5'h5 == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_387 = _T_386 ? _T_45 : _T_385; // @[Mux.scala 80:57]
  wire  _T_388 = 5'h6 == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_389 = _T_388 ? _T_53 : _T_387; // @[Mux.scala 80:57]
  wire  _T_390 = 5'h7 == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_391 = _T_390 ? _T_61 : _T_389; // @[Mux.scala 80:57]
  wire  _T_392 = 5'h8 == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_393 = _T_392 ? _T_69 : _T_391; // @[Mux.scala 80:57]
  wire  _T_394 = 5'h9 == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_395 = _T_394 ? _T_77 : _T_393; // @[Mux.scala 80:57]
  wire  _T_396 = 5'ha == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_397 = _T_396 ? _T_85 : _T_395; // @[Mux.scala 80:57]
  wire  _T_398 = 5'hb == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_399 = _T_398 ? _T_93 : _T_397; // @[Mux.scala 80:57]
  wire  _T_400 = 5'hc == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_401 = _T_400 ? _T_101 : _T_399; // @[Mux.scala 80:57]
  wire  _T_402 = 5'hd == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_403 = _T_402 ? _T_109 : _T_401; // @[Mux.scala 80:57]
  wire  _T_404 = 5'he == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_405 = _T_404 ? _T_117 : _T_403; // @[Mux.scala 80:57]
  wire  _T_406 = 5'hf == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_407 = _T_406 ? _T_125 : _T_405; // @[Mux.scala 80:57]
  wire  _T_408 = 5'h10 == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_409 = _T_408 ? _T_133 : _T_407; // @[Mux.scala 80:57]
  wire  _T_410 = 5'h11 == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_411 = _T_410 ? _T_141 : _T_409; // @[Mux.scala 80:57]
  wire  _T_412 = 5'h12 == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_413 = _T_412 ? _T_149 : _T_411; // @[Mux.scala 80:57]
  wire  _T_414 = 5'h13 == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_415 = _T_414 ? _T_157 : _T_413; // @[Mux.scala 80:57]
  wire  _T_416 = 5'h14 == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_417 = _T_416 ? _T_165 : _T_415; // @[Mux.scala 80:57]
  wire  _T_418 = 5'h15 == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_419 = _T_418 ? _T_173 : _T_417; // @[Mux.scala 80:57]
  wire  _T_420 = 5'h16 == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_421 = _T_420 ? _T_181 : _T_419; // @[Mux.scala 80:57]
  wire  _T_422 = 5'h17 == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_423 = _T_422 ? _T_189 : _T_421; // @[Mux.scala 80:57]
  wire  _T_424 = 5'h18 == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_425 = _T_424 ? _T_197 : _T_423; // @[Mux.scala 80:57]
  wire  _T_426 = 5'h19 == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_427 = _T_426 ? _T_205 : _T_425; // @[Mux.scala 80:57]
  wire  _T_428 = 5'h1a == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_429 = _T_428 ? _T_213 : _T_427; // @[Mux.scala 80:57]
  wire  _T_430 = 5'h1b == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_431 = _T_430 ? _T_221 : _T_429; // @[Mux.scala 80:57]
  wire  _T_432 = 5'h1c == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_433 = _T_432 ? _T_229 : _T_431; // @[Mux.scala 80:57]
  wire  _T_434 = 5'h1d == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_435 = _T_434 ? _T_237 : _T_433; // @[Mux.scala 80:57]
  wire  _T_436 = 5'h1e == io_rdID; // @[Mux.scala 80:60]
  wire [63:0] _T_437 = _T_436 ? _T_245 : _T_435; // @[Mux.scala 80:57]
  wire  _T_438 = 5'h1f == io_rdID; // @[Mux.scala 80:60]
  wire  _T_443 = io_we & _T_3; // @[regFile.scala 68:43]
  reg [63:0] _T_444; // @[Reg.scala 27:20]
  DPIC_RegRead DPIC_RegRead_ins ( // @[regFile.scala 30:33]
    .inst_0(DPIC_RegRead_ins_inst_0),
    .inst_1(DPIC_RegRead_ins_inst_1),
    .inst_2(DPIC_RegRead_ins_inst_2),
    .inst_3(DPIC_RegRead_ins_inst_3),
    .inst_4(DPIC_RegRead_ins_inst_4),
    .inst_5(DPIC_RegRead_ins_inst_5),
    .inst_6(DPIC_RegRead_ins_inst_6),
    .inst_7(DPIC_RegRead_ins_inst_7),
    .inst_8(DPIC_RegRead_ins_inst_8),
    .inst_9(DPIC_RegRead_ins_inst_9),
    .inst_10(DPIC_RegRead_ins_inst_10),
    .inst_11(DPIC_RegRead_ins_inst_11),
    .inst_12(DPIC_RegRead_ins_inst_12),
    .inst_13(DPIC_RegRead_ins_inst_13),
    .inst_14(DPIC_RegRead_ins_inst_14),
    .inst_15(DPIC_RegRead_ins_inst_15),
    .inst_16(DPIC_RegRead_ins_inst_16),
    .inst_17(DPIC_RegRead_ins_inst_17),
    .inst_18(DPIC_RegRead_ins_inst_18),
    .inst_19(DPIC_RegRead_ins_inst_19),
    .inst_20(DPIC_RegRead_ins_inst_20),
    .inst_21(DPIC_RegRead_ins_inst_21),
    .inst_22(DPIC_RegRead_ins_inst_22),
    .inst_23(DPIC_RegRead_ins_inst_23),
    .inst_24(DPIC_RegRead_ins_inst_24),
    .inst_25(DPIC_RegRead_ins_inst_25),
    .inst_26(DPIC_RegRead_ins_inst_26),
    .inst_27(DPIC_RegRead_ins_inst_27),
    .inst_28(DPIC_RegRead_ins_inst_28),
    .inst_29(DPIC_RegRead_ins_inst_29),
    .inst_30(DPIC_RegRead_ins_inst_30),
    .inst_31(DPIC_RegRead_ins_inst_31),
    .pc(DPIC_RegRead_ins_pc)
  );
  assign io_dout1 = _T_314 ? _T_253 : _T_313; // @[regFile.scala 64:12]
  assign io_dout2 = _T_376 ? _T_253 : _T_375; // @[regFile.scala 65:12]
  assign io_rdDout = _T_438 ? _T_253 : _T_437; // @[regFile.scala 66:13]
  assign io_doutWB = _T_444; // @[regFile.scala 68:13]
  assign DPIC_RegRead_ins_inst_0 = 64'h0; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_1 = _T_13; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_2 = _T_21; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_3 = _T_29; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_4 = _T_37; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_5 = _T_45; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_6 = _T_53; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_7 = _T_61; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_8 = _T_69; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_9 = _T_77; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_10 = _T_85; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_11 = _T_93; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_12 = _T_101; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_13 = _T_109; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_14 = _T_117; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_15 = _T_125; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_16 = _T_133; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_17 = _T_141; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_18 = _T_149; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_19 = _T_157; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_20 = _T_165; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_21 = _T_173; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_22 = _T_181; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_23 = _T_189; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_24 = _T_197; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_25 = _T_205; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_26 = _T_213; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_27 = _T_221; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_28 = _T_229; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_29 = _T_237; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_30 = _T_245; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_inst_31 = _T_253; // @[regFile.scala 59:35]
  assign DPIC_RegRead_ins_pc = {{32'd0}, io_pc}; // @[regFile.scala 31:55]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_13 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  _T_21 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  _T_29 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  _T_37 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  _T_45 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  _T_53 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  _T_61 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  _T_69 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  _T_77 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  _T_85 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  _T_93 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  _T_101 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  _T_109 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  _T_117 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  _T_125 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  _T_133 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  _T_141 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  _T_149 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  _T_157 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  _T_165 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  _T_173 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  _T_181 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  _T_189 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  _T_197 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  _T_205 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  _T_213 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  _T_221 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  _T_229 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  _T_237 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  _T_245 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  _T_253 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  _T_444 = _RAND_31[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_12) begin
      _T_13 <= io_din;
    end
    if (_T_20) begin
      _T_21 <= io_din;
    end
    if (_T_28) begin
      _T_29 <= io_din;
    end
    if (_T_36) begin
      _T_37 <= io_din;
    end
    if (_T_44) begin
      _T_45 <= io_din;
    end
    if (_T_52) begin
      _T_53 <= io_din;
    end
    if (_T_60) begin
      _T_61 <= io_din;
    end
    if (_T_68) begin
      _T_69 <= io_din;
    end
    if (_T_76) begin
      _T_77 <= io_din;
    end
    if (_T_84) begin
      _T_85 <= io_din;
    end
    if (_T_92) begin
      _T_93 <= io_din;
    end
    if (_T_100) begin
      _T_101 <= io_din;
    end
    if (_T_108) begin
      _T_109 <= io_din;
    end
    if (_T_116) begin
      _T_117 <= io_din;
    end
    if (_T_124) begin
      _T_125 <= io_din;
    end
    if (_T_132) begin
      _T_133 <= io_din;
    end
    if (_T_140) begin
      _T_141 <= io_din;
    end
    if (_T_148) begin
      _T_149 <= io_din;
    end
    if (_T_156) begin
      _T_157 <= io_din;
    end
    if (_T_164) begin
      _T_165 <= io_din;
    end
    if (_T_172) begin
      _T_173 <= io_din;
    end
    if (_T_180) begin
      _T_181 <= io_din;
    end
    if (_T_188) begin
      _T_189 <= io_din;
    end
    if (_T_196) begin
      _T_197 <= io_din;
    end
    if (_T_204) begin
      _T_205 <= io_din;
    end
    if (_T_212) begin
      _T_213 <= io_din;
    end
    if (_T_220) begin
      _T_221 <= io_din;
    end
    if (_T_228) begin
      _T_229 <= io_din;
    end
    if (_T_236) begin
      _T_237 <= io_din;
    end
    if (_T_244) begin
      _T_245 <= io_din;
    end
    if (_T_252) begin
      _T_253 <= io_din;
    end
    if (reset) begin
      _T_444 <= 64'h0;
    end else if (_T_443) begin
      _T_444 <= io_din;
    end
  end
endmodule
module iDecode(
  input         clock,
  input         reset,
  input  [31:0] io_pc,
  input  [31:0] io_inst,
  input         io_regEn,
  output [63:0] io_dataEx_imme,
  output [63:0] io_dataEx_dOut1,
  output [63:0] io_dataEx_dOut2,
  input  [63:0] io_dataEx_dIn,
  output [63:0] io_dataEx_rdDout,
  output [4:0]  io_rdOut,
  input  [4:0]  io_rdIn,
  output [4:0]  io_rs1,
  output [4:0]  io_rs2,
  output [63:0] io_dOutWB,
  input         blockDMA,
  input         block23,
  input         block1
);
  wire [31:0] imme_io_inst; // @[iDecode.scala 28:19]
  wire [63:0] imme_io_imme; // @[iDecode.scala 28:19]
  wire  rf_clock; // @[iDecode.scala 42:18]
  wire  rf_reset; // @[iDecode.scala 42:18]
  wire [31:0] rf_io_pc; // @[iDecode.scala 42:18]
  wire  rf_io_we; // @[iDecode.scala 42:18]
  wire [4:0] rf_io_rs1; // @[iDecode.scala 42:18]
  wire [4:0] rf_io_rs2; // @[iDecode.scala 42:18]
  wire [4:0] rf_io_rd; // @[iDecode.scala 42:18]
  wire [4:0] rf_io_rdID; // @[iDecode.scala 42:18]
  wire [63:0] rf_io_dout1; // @[iDecode.scala 42:18]
  wire [63:0] rf_io_dout2; // @[iDecode.scala 42:18]
  wire [63:0] rf_io_rdDout; // @[iDecode.scala 42:18]
  wire [63:0] rf_io_din; // @[iDecode.scala 42:18]
  wire [63:0] rf_io_doutWB; // @[iDecode.scala 42:18]
  wire  rf_blockDMA_0; // @[iDecode.scala 42:18]
  wire  rf_block23_0; // @[iDecode.scala 42:18]
  wire  rf_block1_0; // @[iDecode.scala 42:18]
  immeGen imme ( // @[iDecode.scala 28:19]
    .io_inst(imme_io_inst),
    .io_imme(imme_io_imme)
  );
  RF rf ( // @[iDecode.scala 42:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_pc(rf_io_pc),
    .io_we(rf_io_we),
    .io_rs1(rf_io_rs1),
    .io_rs2(rf_io_rs2),
    .io_rd(rf_io_rd),
    .io_rdID(rf_io_rdID),
    .io_dout1(rf_io_dout1),
    .io_dout2(rf_io_dout2),
    .io_rdDout(rf_io_rdDout),
    .io_din(rf_io_din),
    .io_doutWB(rf_io_doutWB),
    .blockDMA_0(rf_blockDMA_0),
    .block23_0(rf_block23_0),
    .block1_0(rf_block1_0)
  );
  assign io_dataEx_imme = imme_io_imme; // @[iDecode.scala 30:18]
  assign io_dataEx_dOut1 = rf_io_dout1; // @[iDecode.scala 48:19]
  assign io_dataEx_dOut2 = rf_io_dout2; // @[iDecode.scala 49:19]
  assign io_dataEx_rdDout = rf_io_rdDout; // @[iDecode.scala 51:20]
  assign io_rdOut = io_inst[11:7]; // @[iDecode.scala 37:12]
  assign io_rs1 = io_inst[19:15]; // @[iDecode.scala 38:10]
  assign io_rs2 = io_inst[24:20]; // @[iDecode.scala 39:10]
  assign io_dOutWB = rf_io_doutWB; // @[iDecode.scala 56:13]
  assign imme_io_inst = io_inst; // @[iDecode.scala 29:16]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_pc = io_pc; // @[iDecode.scala 53:12]
  assign rf_io_we = io_regEn; // @[iDecode.scala 46:12]
  assign rf_io_rs1 = io_inst[19:15]; // @[iDecode.scala 43:13]
  assign rf_io_rs2 = io_inst[24:20]; // @[iDecode.scala 44:13]
  assign rf_io_rd = io_rdIn; // @[iDecode.scala 45:12]
  assign rf_io_rdID = io_inst[11:7]; // @[iDecode.scala 50:14]
  assign rf_io_din = io_dataEx_dIn; // @[iDecode.scala 47:13]
  assign rf_blockDMA_0 = blockDMA;
  assign rf_block23_0 = block23;
  assign rf_block1_0 = block1;
endmodule
module add(
  input         io_cin,
  input  [63:0] io_a,
  input  [63:0] io_b,
  output [63:0] io_sum,
  output        io_cout
);
  wire [64:0] _T_1 = {1'h0,io_a}; // @[Cat.scala 29:58]
  wire [64:0] _T_2 = {1'h0,io_b}; // @[Cat.scala 29:58]
  wire [64:0] _T_4 = _T_1 + _T_2; // @[add.scala 18:31]
  wire [64:0] _GEN_0 = {{64'd0}, io_cin}; // @[add.scala 18:52]
  wire [64:0] _T_6 = _T_4 + _GEN_0; // @[add.scala 18:52]
  assign io_sum = _T_6[63:0]; // @[add.scala 19:12]
  assign io_cout = _T_6[64]; // @[add.scala 20:13]
endmodule
module divR2(
  input         clock,
  input         reset,
  input  [63:0] io_dividend,
  input  [63:0] io_divisor,
  input         io_div_valid,
  input         io_divw,
  input         io_div_signed,
  output        io_out_valid,
  output [63:0] io_quotient,
  output [63:0] io_remainder,
  input         io_block
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  _T_1 = io_dividend[63] & io_div_signed; // @[divR2.scala 22:51]
  wire [63:0] _T_2 = ~io_dividend; // @[divR2.scala 22:70]
  wire [63:0] _T_4 = _T_2 + 64'h1; // @[divR2.scala 22:91]
  wire [63:0] dividend64Real = _T_1 ? _T_4 : io_dividend; // @[divR2.scala 22:27]
  wire  _T_6 = io_divisor[63] & io_div_signed; // @[divR2.scala 23:49]
  wire [63:0] _T_7 = ~io_divisor; // @[divR2.scala 23:68]
  wire [63:0] _T_9 = _T_7 + 64'h1; // @[divR2.scala 23:88]
  wire [63:0] divisor64Real = _T_6 ? _T_9 : io_divisor; // @[divR2.scala 23:26]
  wire  _T_12 = io_dividend[63] ^ io_divisor[63]; // @[divR2.scala 24:42]
  wire  quoSgn64 = _T_12 & io_div_signed; // @[divR2.scala 24:67]
  wire  _T_15 = io_dividend[31] & io_div_signed; // @[divR2.scala 27:48]
  wire [31:0] _T_17 = ~io_dividend[31:0]; // @[divR2.scala 27:67]
  wire [31:0] _T_19 = _T_17 + 32'h1; // @[divR2.scala 27:94]
  wire [31:0] dividend32Real = _T_15 ? _T_19 : io_dividend[31:0]; // @[divR2.scala 27:27]
  wire  _T_22 = io_divisor[31] & io_div_signed; // @[divR2.scala 28:46]
  wire [31:0] _T_24 = ~io_divisor[31:0]; // @[divR2.scala 28:65]
  wire [31:0] _T_26 = _T_24 + 32'h1; // @[divR2.scala 28:91]
  wire [31:0] divisor32Real = _T_22 ? _T_26 : io_divisor[31:0]; // @[divR2.scala 28:26]
  wire  _T_30 = io_dividend[31] ^ io_divisor[31]; // @[divR2.scala 29:39]
  wire  quoSgn32 = _T_30 & io_div_signed; // @[divR2.scala 29:61]
  reg [1:0] stateReg; // @[divR2.scala 36:25]
  wire  isDiv32 = stateReg == 2'h1; // @[divR2.scala 38:25]
  wire  isDiv64 = stateReg == 2'h2; // @[divR2.scala 39:26]
  reg [5:0] cnt; // @[divR2.scala 41:20]
  wire [1:0] _T_32 = {io_div_valid,io_divw}; // @[Cat.scala 29:58]
  wire  _T_33 = 2'h3 == _T_32; // @[Mux.scala 80:60]
  wire  _T_35 = 2'h2 == _T_32; // @[Mux.scala 80:60]
  wire  _T_36 = cnt == 6'h1f; // @[divR2.scala 50:26]
  wire  _T_37 = cnt == 6'h3f; // @[divR2.scala 51:26]
  wire  _T_38 = 2'h1 == stateReg; // @[Mux.scala 80:60]
  wire  _T_40 = 2'h2 == stateReg; // @[Mux.scala 80:60]
  wire  _T_42 = 2'h3 == stateReg; // @[Mux.scala 80:60]
  wire  _T_44 = isDiv32 | isDiv64; // @[divR2.scala 64:21]
  wire [5:0] _T_46 = cnt + 6'h1; // @[divR2.scala 64:38]
  reg [127:0] dividendReg; // @[divR2.scala 67:28]
  reg [63:0] resReg; // @[divR2.scala 68:23]
  wire [127:0] _T_51 = {96'h0,dividend32Real}; // @[Cat.scala 29:58]
  wire [127:0] _T_52 = {64'h0,dividend64Real}; // @[Cat.scala 29:58]
  wire [32:0] subed32 = dividendReg[63:31]; // @[divR2.scala 96:27]
  wire [32:0] _GEN_0 = {{1'd0}, divisor32Real}; // @[divR2.scala 97:26]
  wire [32:0] subRes32 = subed32 - _GEN_0; // @[divR2.scala 97:26]
  wire [31:0] rem32M = subRes32[32] ? subed32[31:0] : subRes32[31:0]; // @[divR2.scala 98:16]
  wire [127:0] div32DividendMux = {64'h0,rem32M,dividendReg[30:0],1'h0}; // @[Cat.scala 29:58]
  wire [64:0] subed64 = dividendReg[127:63]; // @[divR2.scala 92:29]
  wire [64:0] _GEN_1 = {{1'd0}, divisor64Real}; // @[divR2.scala 93:26]
  wire [64:0] subRes64 = subed64 - _GEN_1; // @[divR2.scala 93:26]
  wire [63:0] rem64M = subRes64[64] ? subed64[63:0] : subRes64[63:0]; // @[divR2.scala 94:16]
  wire [127:0] div64DividendMux = {rem64M,dividendReg[62:0],1'h0}; // @[Cat.scala 29:58]
  wire  _T_79 = ~subRes32[32]; // @[divR2.scala 105:38]
  wire [63:0] _T_80 = {resReg[62:0],_T_79}; // @[Cat.scala 29:58]
  wire  _T_83 = ~subRes64[64]; // @[divR2.scala 106:38]
  wire [63:0] _T_84 = {resReg[62:0],_T_83}; // @[Cat.scala 29:58]
  wire [63:0] _T_91 = ~resReg; // @[divR2.scala 111:35]
  wire [63:0] _T_93 = _T_91 + 64'h1; // @[divR2.scala 111:53]
  wire [63:0] res64Out = quoSgn64 ? _T_93 : resReg; // @[divR2.scala 111:21]
  wire [63:0] _T_95 = ~dividendReg[127:64]; // @[divR2.scala 112:32]
  wire [63:0] _T_97 = _T_95 + 64'h1; // @[divR2.scala 112:63]
  wire [63:0] rem64Out = _T_1 ? _T_97 : dividendReg[127:64]; // @[divR2.scala 112:20]
  wire [31:0] _T_101 = ~resReg[31:0]; // @[divR2.scala 114:56]
  wire [31:0] _T_103 = _T_101 + 32'h1; // @[divR2.scala 114:79]
  wire [63:0] _T_104 = {32'hffffffff,_T_103}; // @[Cat.scala 29:58]
  wire [63:0] res32out = quoSgn32 ? _T_104 : resReg; // @[divR2.scala 114:21]
  wire [31:0] _T_107 = ~dividendReg[63:32]; // @[divR2.scala 116:56]
  wire [31:0] _T_109 = _T_107 + 32'h1; // @[divR2.scala 116:85]
  wire [63:0] _T_110 = {32'hffffffff,_T_109}; // @[Cat.scala 29:58]
  wire [63:0] _T_113 = {32'h0,dividendReg[63:32]}; // @[Cat.scala 29:58]
  wire [63:0] rem32Out = _T_15 ? _T_110 : _T_113; // @[divR2.scala 116:21]
  assign io_out_valid = stateReg == 2'h3; // @[divR2.scala 124:16]
  assign io_quotient = io_divw ? res32out : res64Out; // @[divR2.scala 120:15]
  assign io_remainder = io_divw ? rem32Out : rem64Out; // @[divR2.scala 121:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  cnt = _RAND_1[5:0];
  _RAND_2 = {4{`RANDOM}};
  dividendReg = _RAND_2[127:0];
  _RAND_3 = {2{`RANDOM}};
  resReg = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      stateReg <= 2'h0;
    end else if (_T_42) begin
      if (io_block) begin
        stateReg <= 2'h3;
      end else begin
        stateReg <= 2'h0;
      end
    end else if (_T_40) begin
      if (_T_37) begin
        stateReg <= 2'h3;
      end else begin
        stateReg <= 2'h2;
      end
    end else if (_T_38) begin
      if (_T_36) begin
        stateReg <= 2'h3;
      end else begin
        stateReg <= 2'h1;
      end
    end else if (_T_35) begin
      stateReg <= 2'h2;
    end else if (_T_33) begin
      stateReg <= 2'h1;
    end else begin
      stateReg <= 2'h0;
    end
    if (reset) begin
      cnt <= 6'h0;
    end else if (_T_44) begin
      cnt <= _T_46;
    end else begin
      cnt <= 6'h0;
    end
    if (reset) begin
      dividendReg <= 128'h0;
    end else if (!(_T_42)) begin
      if (_T_40) begin
        dividendReg <= div64DividendMux;
      end else if (_T_38) begin
        dividendReg <= div32DividendMux;
      end else if (_T_35) begin
        dividendReg <= _T_52;
      end else if (_T_33) begin
        dividendReg <= _T_51;
      end else begin
        dividendReg <= 128'h0;
      end
    end
    if (reset) begin
      resReg <= 64'h0;
    end else if (!(_T_42)) begin
      if (_T_40) begin
        resReg <= _T_84;
      end else if (_T_38) begin
        resReg <= _T_80;
      end else begin
        resReg <= 64'h0;
      end
    end
  end
endmodule
module mul(
  input         clock,
  input         reset,
  input         io_mul_valid,
  input  [63:0] io_multiplicand,
  input  [63:0] io_multiplier,
  output        io_out_valid,
  output [63:0] io_result_low,
  input         io_block
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [127:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] _T; // @[mul.scala 43:27]
  wire  _T_1 = _T == 2'h0; // @[mul.scala 44:27]
  wire  _T_2 = _T == 2'h1; // @[mul.scala 45:26]
  wire  _T_6 = 2'h0 == _T; // @[Mux.scala 80:60]
  wire  _T_8 = 2'h1 == _T; // @[Mux.scala 80:60]
  wire  _T_10 = 2'h2 == _T; // @[Mux.scala 80:60]
  wire  _T_12 = _T_1 & io_mul_valid; // @[mul.scala 59:64]
  reg [63:0] _T_13; // @[Reg.scala 27:20]
  reg [63:0] _T_15; // @[Reg.scala 27:20]
  wire [127:0] _T_16 = _T_13 * _T_15; // @[mul.scala 61:31]
  reg [127:0] _T_17; // @[Reg.scala 27:20]
  assign io_out_valid = _T == 2'h2; // @[mul.scala 66:18]
  assign io_result_low = _T_17[63:0]; // @[mul.scala 64:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  _T_13 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  _T_15 = _RAND_2[63:0];
  _RAND_3 = {4{`RANDOM}};
  _T_17 = _RAND_3[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T <= 2'h0;
    end else if (_T_10) begin
      if (io_block) begin
        _T <= 2'h2;
      end else begin
        _T <= 2'h0;
      end
    end else if (_T_8) begin
      _T <= 2'h2;
    end else if (_T_6) begin
      if (io_mul_valid) begin
        _T <= 2'h1;
      end else begin
        _T <= 2'h0;
      end
    end else begin
      _T <= 2'h0;
    end
    if (reset) begin
      _T_13 <= 64'h0;
    end else if (_T_12) begin
      _T_13 <= io_multiplicand;
    end
    if (reset) begin
      _T_15 <= 64'h0;
    end else if (_T_12) begin
      _T_15 <= io_multiplier;
    end
    if (reset) begin
      _T_17 <= 128'h0;
    end else if (_T_2) begin
      _T_17 <= _T_16;
    end
  end
endmodule
module ALU(
  input         clock,
  input         reset,
  input  [63:0] io_srcA,
  input  [63:0] io_srcB,
  input  [4:0]  io_ALUCtrl,
  output [63:0] io_ALUResult,
  input         block23_0,
  output        block1_0
);
  wire  addIns_io_cin; // @[ALU.scala 22:22]
  wire [63:0] addIns_io_a; // @[ALU.scala 22:22]
  wire [63:0] addIns_io_b; // @[ALU.scala 22:22]
  wire [63:0] addIns_io_sum; // @[ALU.scala 22:22]
  wire  addIns_io_cout; // @[ALU.scala 22:22]
  wire  divR2Ins_clock; // @[ALU.scala 31:23]
  wire  divR2Ins_reset; // @[ALU.scala 31:23]
  wire [63:0] divR2Ins_io_dividend; // @[ALU.scala 31:23]
  wire [63:0] divR2Ins_io_divisor; // @[ALU.scala 31:23]
  wire  divR2Ins_io_div_valid; // @[ALU.scala 31:23]
  wire  divR2Ins_io_divw; // @[ALU.scala 31:23]
  wire  divR2Ins_io_div_signed; // @[ALU.scala 31:23]
  wire  divR2Ins_io_out_valid; // @[ALU.scala 31:23]
  wire [63:0] divR2Ins_io_quotient; // @[ALU.scala 31:23]
  wire [63:0] divR2Ins_io_remainder; // @[ALU.scala 31:23]
  wire  divR2Ins_io_block; // @[ALU.scala 31:23]
  wire  mulIns_clock; // @[ALU.scala 46:22]
  wire  mulIns_reset; // @[ALU.scala 46:22]
  wire  mulIns_io_mul_valid; // @[ALU.scala 46:22]
  wire [63:0] mulIns_io_multiplicand; // @[ALU.scala 46:22]
  wire [63:0] mulIns_io_multiplier; // @[ALU.scala 46:22]
  wire  mulIns_io_out_valid; // @[ALU.scala 46:22]
  wire [63:0] mulIns_io_result_low; // @[ALU.scala 46:22]
  wire  mulIns_io_block; // @[ALU.scala 46:22]
  wire  _T = io_ALUCtrl == 5'h1; // @[ALU.scala 24:69]
  wire  _T_2 = io_ALUCtrl == 5'h5; // @[ALU.scala 24:69]
  wire  _T_3 = _T | _T_2; // @[ALU.scala 24:56]
  wire  _T_4 = io_ALUCtrl == 5'h10; // @[ALU.scala 24:69]
  wire  _T_5 = _T_3 | _T_4; // @[ALU.scala 24:56]
  wire  _T_7 = _T_5 | _T_2; // @[ALU.scala 24:56]
  wire  _T_8 = io_ALUCtrl == 5'h7; // @[ALU.scala 24:69]
  wire  _T_9 = _T_7 | _T_8; // @[ALU.scala 24:56]
  wire  _T_10 = io_ALUCtrl == 5'h1b; // @[ALU.scala 24:69]
  wire  _T_11 = _T_9 | _T_10; // @[ALU.scala 24:56]
  wire  _T_12 = io_ALUCtrl == 5'h1c; // @[ALU.scala 24:69]
  wire  sub = _T_11 | _T_12; // @[ALU.scala 24:56]
  wire [63:0] srcBInv = ~io_srcB; // @[ALU.scala 25:18]
  wire  _T_14 = io_ALUCtrl == 5'h11; // @[ALU.scala 33:79]
  wire  _T_16 = io_ALUCtrl == 5'h12; // @[ALU.scala 33:79]
  wire  _T_17 = _T_14 | _T_16; // @[ALU.scala 33:66]
  wire  _T_18 = io_ALUCtrl == 5'h14; // @[ALU.scala 33:79]
  wire  _T_19 = _T_17 | _T_18; // @[ALU.scala 33:66]
  wire  _T_20 = io_ALUCtrl == 5'h15; // @[ALU.scala 33:79]
  wire  _T_21 = _T_19 | _T_20; // @[ALU.scala 33:66]
  wire  _T_22 = io_ALUCtrl == 5'h17; // @[ALU.scala 33:79]
  wire  _T_23 = _T_21 | _T_22; // @[ALU.scala 33:66]
  wire  _T_24 = io_ALUCtrl == 5'h18; // @[ALU.scala 33:79]
  wire  _T_25 = _T_23 | _T_24; // @[ALU.scala 33:66]
  wire  _T_26 = io_ALUCtrl == 5'h19; // @[ALU.scala 33:79]
  wire  _T_27 = _T_25 | _T_26; // @[ALU.scala 33:66]
  wire  _T_28 = io_ALUCtrl == 5'h1d; // @[ALU.scala 33:79]
  wire  _T_39 = _T_18 | _T_20; // @[ALU.scala 37:68]
  wire  _T_41 = _T_39 | _T_24; // @[ALU.scala 37:68]
  wire [63:0] srcAUSignW = {32'h0,io_srcA[31:0]}; // @[Cat.scala 29:58]
  wire [63:0] srcBUSignW = {32'h0,io_srcB[31:0]}; // @[Cat.scala 29:58]
  wire  _T_45 = io_ALUCtrl == 5'h13; // @[ALU.scala 50:79]
  wire  _T_47 = io_ALUCtrl == 5'h16; // @[ALU.scala 50:79]
  wire [5:0] shamt = io_srcB[5:0]; // @[ALU.scala 61:22]
  wire [63:0] _T_53 = $signed(io_srcA) >>> shamt; // @[ALU.scala 65:42]
  wire [63:0] _T_54 = io_srcA >> shamt; // @[ALU.scala 66:25]
  wire [126:0] _GEN_0 = {{63'd0}, io_srcA}; // @[ALU.scala 67:25]
  wire [126:0] _T_55 = _GEN_0 << shamt; // @[ALU.scala 67:25]
  wire  _T_57 = ~addIns_io_cout; // @[ALU.scala 69:16]
  wire [63:0] _T_58 = io_srcA & io_srcB; // @[ALU.scala 70:25]
  wire [63:0] _T_59 = io_srcA | io_srcB; // @[ALU.scala 71:24]
  wire [63:0] _T_60 = io_srcA ^ io_srcB; // @[ALU.scala 72:25]
  wire  _T_61 = io_srcA != io_srcB; // @[ALU.scala 73:32]
  wire [63:0] _T_62 = {63'h0,_T_61}; // @[Cat.scala 29:58]
  wire [31:0] _T_64 = io_srcA[31:0] >> shamt; // @[ALU.scala 74:48]
  wire [31:0] _T_67 = _T_64[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_68 = {_T_67,_T_64}; // @[Cat.scala 29:58]
  wire [31:0] _T_72 = addIns_io_sum[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_73 = {_T_72,addIns_io_sum[31:0]}; // @[Cat.scala 29:58]
  wire [94:0] _GEN_1 = {{63'd0}, io_srcA[31:0]}; // @[ALU.scala 76:48]
  wire [94:0] _T_75 = _GEN_1 << shamt; // @[ALU.scala 76:48]
  wire [31:0] _T_79 = _T_75[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_80 = {_T_79,_T_75[31:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_82 = io_srcA[31:0]; // @[ALU.scala 77:41]
  wire [31:0] _T_84 = $signed(_T_82) >>> shamt; // @[ALU.scala 77:65]
  wire [31:0] _T_87 = _T_84[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_88 = {_T_87,_T_84}; // @[Cat.scala 29:58]
  wire [31:0] _T_97 = divR2Ins_io_quotient[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_98 = {_T_97,divR2Ins_io_quotient[31:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_102 = divR2Ins_io_remainder[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_103 = {_T_102,divR2Ins_io_remainder[31:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_107 = mulIns_io_result_low[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_108 = {_T_107,mulIns_io_result_low[31:0]}; // @[Cat.scala 29:58]
  wire  _T_119 = io_srcA == io_srcB; // @[ALU.scala 88:24]
  wire  _T_121 = ~addIns_io_sum[63]; // @[ALU.scala 91:16]
  wire  _T_122 = 5'h0 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [63:0] _T_123 = _T_122 ? addIns_io_sum : 64'h0; // @[Mux.scala 80:57]
  wire  _T_124 = 5'h1 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [63:0] _T_125 = _T_124 ? addIns_io_sum : _T_123; // @[Mux.scala 80:57]
  wire  _T_126 = 5'h9 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [63:0] _T_127 = _T_126 ? _T_53 : _T_125; // @[Mux.scala 80:57]
  wire  _T_128 = 5'h8 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [63:0] _T_129 = _T_128 ? _T_54 : _T_127; // @[Mux.scala 80:57]
  wire  _T_130 = 5'h6 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_131 = _T_130 ? _T_55 : {{63'd0}, _T_129}; // @[Mux.scala 80:57]
  wire  _T_132 = 5'h5 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_133 = _T_132 ? {{126'd0}, addIns_io_sum[63]} : _T_131; // @[Mux.scala 80:57]
  wire  _T_134 = 5'h7 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_135 = _T_134 ? {{126'd0}, _T_57} : _T_133; // @[Mux.scala 80:57]
  wire  _T_136 = 5'h2 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_137 = _T_136 ? {{63'd0}, _T_58} : _T_135; // @[Mux.scala 80:57]
  wire  _T_138 = 5'h3 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_139 = _T_138 ? {{63'd0}, _T_59} : _T_137; // @[Mux.scala 80:57]
  wire  _T_140 = 5'h4 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_141 = _T_140 ? {{63'd0}, _T_60} : _T_139; // @[Mux.scala 80:57]
  wire  _T_142 = 5'hb == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_143 = _T_142 ? {{63'd0}, _T_62} : _T_141; // @[Mux.scala 80:57]
  wire  _T_144 = 5'hc == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_145 = _T_144 ? {{63'd0}, _T_68} : _T_143; // @[Mux.scala 80:57]
  wire  _T_146 = 5'hd == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_147 = _T_146 ? {{63'd0}, _T_73} : _T_145; // @[Mux.scala 80:57]
  wire  _T_148 = 5'he == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_149 = _T_148 ? {{63'd0}, _T_80} : _T_147; // @[Mux.scala 80:57]
  wire  _T_150 = 5'hf == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_151 = _T_150 ? {{63'd0}, _T_88} : _T_149; // @[Mux.scala 80:57]
  wire  _T_152 = 5'h10 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_153 = _T_152 ? {{63'd0}, _T_73} : _T_151; // @[Mux.scala 80:57]
  wire  _T_154 = 5'h11 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_155 = _T_154 ? {{63'd0}, _T_98} : _T_153; // @[Mux.scala 80:57]
  wire  _T_156 = 5'h12 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_157 = _T_156 ? {{63'd0}, _T_103} : _T_155; // @[Mux.scala 80:57]
  wire  _T_158 = 5'h13 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_159 = _T_158 ? {{63'd0}, _T_108} : _T_157; // @[Mux.scala 80:57]
  wire  _T_160 = 5'h14 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_161 = _T_160 ? {{63'd0}, _T_103} : _T_159; // @[Mux.scala 80:57]
  wire  _T_162 = 5'h15 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_163 = _T_162 ? {{63'd0}, _T_98} : _T_161; // @[Mux.scala 80:57]
  wire  _T_164 = 5'h16 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_165 = _T_164 ? {{63'd0}, mulIns_io_result_low} : _T_163; // @[Mux.scala 80:57]
  wire  _T_166 = 5'h17 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_167 = _T_166 ? {{63'd0}, divR2Ins_io_quotient} : _T_165; // @[Mux.scala 80:57]
  wire  _T_168 = 5'h18 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_169 = _T_168 ? {{63'd0}, divR2Ins_io_remainder} : _T_167; // @[Mux.scala 80:57]
  wire  _T_170 = 5'h19 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_171 = _T_170 ? {{63'd0}, divR2Ins_io_quotient} : _T_169; // @[Mux.scala 80:57]
  wire  _T_172 = 5'h1a == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_173 = _T_172 ? {{126'd0}, _T_119} : _T_171; // @[Mux.scala 80:57]
  wire  _T_174 = 5'h1b == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_175 = _T_174 ? {{126'd0}, addIns_io_cout} : _T_173; // @[Mux.scala 80:57]
  wire  _T_176 = 5'h1c == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_177 = _T_176 ? {{126'd0}, _T_121} : _T_175; // @[Mux.scala 80:57]
  wire  _T_178 = 5'h1d == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_179 = _T_178 ? {{63'd0}, divR2Ins_io_remainder} : _T_177; // @[Mux.scala 80:57]
  wire  _T_180 = 5'ha == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_181 = _T_180 ? {{63'd0}, io_srcA} : _T_179; // @[Mux.scala 80:57]
  wire  _T_182 = ~divR2Ins_io_out_valid; // @[ALU.scala 98:38]
  wire  _T_183 = divR2Ins_io_div_valid & _T_182; // @[ALU.scala 98:35]
  wire  _T_184 = ~mulIns_io_out_valid; // @[ALU.scala 98:87]
  wire  _T_185 = mulIns_io_mul_valid & _T_184; // @[ALU.scala 98:84]
  wire  _T_186 = _T_183 | _T_185; // @[ALU.scala 98:61]
  wire  block1 = _T_186; // @[ALU.scala 97:20 ALU.scala 98:10]
  add addIns ( // @[ALU.scala 22:22]
    .io_cin(addIns_io_cin),
    .io_a(addIns_io_a),
    .io_b(addIns_io_b),
    .io_sum(addIns_io_sum),
    .io_cout(addIns_io_cout)
  );
  divR2 divR2Ins ( // @[ALU.scala 31:23]
    .clock(divR2Ins_clock),
    .reset(divR2Ins_reset),
    .io_dividend(divR2Ins_io_dividend),
    .io_divisor(divR2Ins_io_divisor),
    .io_div_valid(divR2Ins_io_div_valid),
    .io_divw(divR2Ins_io_divw),
    .io_div_signed(divR2Ins_io_div_signed),
    .io_out_valid(divR2Ins_io_out_valid),
    .io_quotient(divR2Ins_io_quotient),
    .io_remainder(divR2Ins_io_remainder),
    .io_block(divR2Ins_io_block)
  );
  mul mulIns ( // @[ALU.scala 46:22]
    .clock(mulIns_clock),
    .reset(mulIns_reset),
    .io_mul_valid(mulIns_io_mul_valid),
    .io_multiplicand(mulIns_io_multiplicand),
    .io_multiplier(mulIns_io_multiplier),
    .io_out_valid(mulIns_io_out_valid),
    .io_result_low(mulIns_io_result_low),
    .io_block(mulIns_io_block)
  );
  assign io_ALUResult = _T_181[63:0]; // @[ALU.scala 95:16]
  assign block1_0 = block1;
  assign addIns_io_cin = _T_11 | _T_12; // @[ALU.scala 26:17]
  assign addIns_io_a = io_srcA; // @[ALU.scala 27:15]
  assign addIns_io_b = sub ? srcBInv : io_srcB; // @[ALU.scala 28:55]
  assign divR2Ins_clock = clock;
  assign divR2Ins_reset = reset;
  assign divR2Ins_io_dividend = io_srcA; // @[ALU.scala 38:24]
  assign divR2Ins_io_divisor = io_srcB; // @[ALU.scala 39:23]
  assign divR2Ins_io_div_valid = _T_27 | _T_28; // @[ALU.scala 40:25]
  assign divR2Ins_io_divw = _T_19 | _T_20; // @[ALU.scala 41:20]
  assign divR2Ins_io_div_signed = _T_41 | _T_26; // @[ALU.scala 42:26]
  assign divR2Ins_io_block = block23_0; // @[ALU.scala 111:21]
  assign mulIns_clock = clock;
  assign mulIns_reset = reset;
  assign mulIns_io_mul_valid = _T_45 | _T_47; // @[ALU.scala 55:23]
  assign mulIns_io_multiplicand = _T_45 ? srcAUSignW : io_srcA; // @[ALU.scala 56:26]
  assign mulIns_io_multiplier = _T_45 ? srcBUSignW : io_srcB; // @[ALU.scala 57:24]
  assign mulIns_io_block = block23_0; // @[ALU.scala 110:19]
endmodule
module CSR(
  input         clock,
  input         reset,
  input         io_csrrwen,
  input         io_csrswen,
  input         io_csrrsien,
  input         io_csrrcien,
  input         io_csrrcen,
  input         io_csrrwien,
  input         io_ecall,
  input  [63:0] io_rs1,
  input  [11:0] io_imme,
  input  [63:0] io_pc,
  input  [4:0]  io_uimm,
  output [63:0] io_rd,
  output [63:0] io_mtvec,
  output [63:0] io_mepc,
  input         io_mret,
  input         intrTimeCnt_0,
  output        startTimeCnt_0,
  input         blockDMA_0,
  input         block23_0,
  input         block1_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  _T = io_pc != 64'h0; // @[CSR.scala 37:35]
  wire  intr = intrTimeCnt_0 & _T; // @[CSR.scala 37:26]
  wire  _T_1 = io_csrrwen | io_csrswen; // @[CSR.scala 54:26]
  wire  _T_2 = _T_1 | io_csrrcen; // @[CSR.scala 54:38]
  wire  _T_3 = _T_2 | io_csrrsien; // @[CSR.scala 54:52]
  wire  _T_4 = _T_3 | io_csrrcien; // @[CSR.scala 54:67]
  wire  csren = _T_4 | io_csrrwien; // @[CSR.scala 54:82]
  wire [5:0] sel1H = {io_csrrwien,io_csrrcien,io_csrrsien,io_csrrcen,io_csrswen,io_csrrwen}; // @[Cat.scala 29:58]
  wire [63:0] uimmext = {59'h0,io_uimm}; // @[Cat.scala 29:58]
  wire  _T_9 = io_imme == 12'h341; // @[CSR.scala 58:48]
  wire  _T_10 = csren & _T_9; // @[CSR.scala 58:36]
  wire  _T_11 = io_ecall | _T_10; // @[CSR.scala 58:25]
  wire  mepcen = _T_11 | intr; // @[CSR.scala 58:58]
  wire  _T_12 = io_ecall | intr; // @[CSR.scala 61:14]
  reg [63:0] mepcins; // @[Reg.scala 27:20]
  wire [63:0] _T_13 = io_rs1 | mepcins; // @[CSR.scala 67:15]
  wire [63:0] _T_14 = ~io_rs1; // @[CSR.scala 68:10]
  wire [63:0] _T_15 = _T_14 & mepcins; // @[CSR.scala 68:28]
  wire [63:0] _T_16 = uimmext | mepcins; // @[CSR.scala 69:17]
  wire [63:0] _T_17 = ~uimmext; // @[CSR.scala 70:10]
  wire [63:0] _T_18 = _T_17 & mepcins; // @[CSR.scala 70:29]
  wire [63:0] _T_25 = sel1H[0] ? io_rs1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_26 = sel1H[1] ? _T_13 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_27 = sel1H[2] ? _T_15 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_28 = sel1H[3] ? _T_16 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_29 = sel1H[4] ? _T_18 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_30 = sel1H[5] ? uimmext : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_31 = _T_25 | _T_26; // @[Mux.scala 27:72]
  wire [63:0] _T_32 = _T_31 | _T_27; // @[Mux.scala 27:72]
  wire [63:0] _T_33 = _T_32 | _T_28; // @[Mux.scala 27:72]
  wire [63:0] _T_34 = _T_33 | _T_29; // @[Mux.scala 27:72]
  wire [63:0] _T_35 = _T_34 | _T_30; // @[Mux.scala 27:72]
  wire  _T_37 = block1_0 | block23_0; // @[CSR.scala 75:56]
  wire  _T_38 = _T_37 | blockDMA_0; // @[CSR.scala 75:66]
  wire  _T_39 = ~_T_38; // @[CSR.scala 75:47]
  wire  _T_40 = mepcen & _T_39; // @[CSR.scala 75:44]
  wire  _T_42 = io_imme == 12'h342; // @[CSR.scala 77:49]
  wire  _T_43 = csren & _T_42; // @[CSR.scala 77:37]
  wire  _T_44 = io_ecall | _T_43; // @[CSR.scala 77:27]
  wire  mcauseen = _T_44 | intr; // @[CSR.scala 77:61]
  reg [63:0] mcauseins; // @[Reg.scala 27:20]
  wire [63:0] _T_45 = io_rs1 | mcauseins; // @[CSR.scala 89:16]
  wire [63:0] _T_47 = _T_14 & mcauseins; // @[CSR.scala 90:28]
  wire [63:0] _T_48 = uimmext | mcauseins; // @[CSR.scala 91:17]
  wire [63:0] _T_50 = _T_17 & mcauseins; // @[CSR.scala 92:29]
  wire [63:0] _T_58 = sel1H[1] ? _T_45 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_59 = sel1H[2] ? _T_47 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_60 = sel1H[3] ? _T_48 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_61 = sel1H[4] ? _T_50 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_63 = _T_25 | _T_58; // @[Mux.scala 27:72]
  wire [63:0] _T_64 = _T_63 | _T_59; // @[Mux.scala 27:72]
  wire [63:0] _T_65 = _T_64 | _T_60; // @[Mux.scala 27:72]
  wire [63:0] _T_66 = _T_65 | _T_61; // @[Mux.scala 27:72]
  wire [63:0] _T_67 = _T_66 | _T_30; // @[Mux.scala 27:72]
  wire  _T_73 = mcauseen & _T_39; // @[CSR.scala 97:50]
  wire  _T_75 = io_imme == 12'h305; // @[CSR.scala 99:37]
  wire  mtvecen = csren & _T_75; // @[CSR.scala 99:25]
  reg [63:0] mtvecins; // @[Reg.scala 27:20]
  wire [63:0] _T_76 = io_rs1 | mtvecins; // @[CSR.scala 105:14]
  wire [63:0] _T_78 = _T_14 & mtvecins; // @[CSR.scala 106:26]
  wire [63:0] _T_79 = uimmext | mtvecins; // @[CSR.scala 107:15]
  wire [63:0] _T_81 = _T_17 & mtvecins; // @[CSR.scala 108:27]
  wire [63:0] _T_89 = sel1H[1] ? _T_76 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_90 = sel1H[2] ? _T_78 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_91 = sel1H[3] ? _T_79 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_92 = sel1H[4] ? _T_81 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_94 = _T_25 | _T_89; // @[Mux.scala 27:72]
  wire [63:0] _T_95 = _T_94 | _T_90; // @[Mux.scala 27:72]
  wire [63:0] _T_96 = _T_95 | _T_91; // @[Mux.scala 27:72]
  wire [63:0] _T_97 = _T_96 | _T_92; // @[Mux.scala 27:72]
  wire [63:0] mtvecval = _T_97 | _T_30; // @[Mux.scala 27:72]
  wire  _T_100 = _T_37 | intr; // @[CSR.scala 112:70]
  wire  _T_101 = _T_100 | blockDMA_0; // @[CSR.scala 112:77]
  wire  _T_102 = ~_T_101; // @[CSR.scala 112:50]
  wire  _T_103 = mtvecen & _T_102; // @[CSR.scala 112:47]
  wire  _T_105 = io_imme == 12'h300; // @[CSR.scala 114:40]
  wire  _T_106 = csren & _T_105; // @[CSR.scala 114:28]
  wire  _T_107 = _T_106 | io_ecall; // @[CSR.scala 114:54]
  wire  _T_108 = _T_107 | intr; // @[CSR.scala 114:65]
  wire  mstatusen = _T_108 | io_mret; // @[CSR.scala 114:73]
  reg [63:0] mstatusins; // @[Reg.scala 27:20]
  wire [63:0] _T_117 = {mstatusins[63:8],mstatusins[3],mstatusins[6:4],1'h0,mstatusins[2:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_125 = {mstatusins[63:8],1'h1,mstatusins[6:4],mstatusins[7],mstatusins[2:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_126 = io_rs1 | mstatusins; // @[CSR.scala 127:14]
  wire [63:0] _T_128 = _T_14 & mstatusins; // @[CSR.scala 128:26]
  wire [63:0] _T_129 = uimmext | mstatusins; // @[CSR.scala 129:15]
  wire [63:0] _T_131 = _T_17 & mstatusins; // @[CSR.scala 130:27]
  wire [63:0] _T_139 = sel1H[1] ? _T_126 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_140 = sel1H[2] ? _T_128 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_141 = sel1H[3] ? _T_129 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_142 = sel1H[4] ? _T_131 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_144 = _T_25 | _T_139; // @[Mux.scala 27:72]
  wire [63:0] _T_145 = _T_144 | _T_140; // @[Mux.scala 27:72]
  wire [63:0] _T_146 = _T_145 | _T_141; // @[Mux.scala 27:72]
  wire [63:0] _T_147 = _T_146 | _T_142; // @[Mux.scala 27:72]
  wire [63:0] _T_148 = _T_147 | _T_30; // @[Mux.scala 27:72]
  wire  _T_154 = mstatusen & _T_39; // @[CSR.scala 151:73]
  wire  _T_156 = io_imme == 12'h304; // @[CSR.scala 153:36]
  wire  miecen = csren & _T_156; // @[CSR.scala 153:24]
  reg [63:0] mieins; // @[Reg.scala 27:20]
  wire [63:0] _T_157 = io_rs1 | mieins; // @[CSR.scala 159:14]
  wire [63:0] _T_159 = _T_14 & mieins; // @[CSR.scala 160:26]
  wire [63:0] _T_160 = uimmext | mieins; // @[CSR.scala 161:15]
  wire [63:0] _T_162 = _T_17 & mieins; // @[CSR.scala 162:27]
  wire [63:0] _T_170 = sel1H[1] ? _T_157 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_171 = sel1H[2] ? _T_159 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_172 = sel1H[3] ? _T_160 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_173 = sel1H[4] ? _T_162 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_175 = _T_25 | _T_170; // @[Mux.scala 27:72]
  wire [63:0] _T_176 = _T_175 | _T_171; // @[Mux.scala 27:72]
  wire [63:0] _T_177 = _T_176 | _T_172; // @[Mux.scala 27:72]
  wire [63:0] _T_178 = _T_177 | _T_173; // @[Mux.scala 27:72]
  wire [63:0] mieval = _T_178 | _T_30; // @[Mux.scala 27:72]
  wire  _T_184 = miecen & _T_102; // @[CSR.scala 166:41]
  wire  _T_186 = io_imme == 12'h344; // @[CSR.scala 168:35]
  wire  _T_187 = csren & _T_186; // @[CSR.scala 168:23]
  wire  mipcen = _T_187 | intr; // @[CSR.scala 168:45]
  reg [63:0] mipins; // @[Reg.scala 27:20]
  wire [63:0] _T_191 = {mipins[63:8],1'h1,mipins[6:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_192 = io_rs1 | mipins; // @[CSR.scala 177:14]
  wire [63:0] _T_194 = _T_14 & mipins; // @[CSR.scala 178:26]
  wire [63:0] _T_195 = uimmext | mipins; // @[CSR.scala 179:15]
  wire [63:0] _T_197 = _T_17 & mipins; // @[CSR.scala 180:27]
  wire [63:0] _T_205 = sel1H[1] ? _T_192 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_206 = sel1H[2] ? _T_194 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_207 = sel1H[3] ? _T_195 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_208 = sel1H[4] ? _T_197 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_210 = _T_25 | _T_205; // @[Mux.scala 27:72]
  wire [63:0] _T_211 = _T_210 | _T_206; // @[Mux.scala 27:72]
  wire [63:0] _T_212 = _T_211 | _T_207; // @[Mux.scala 27:72]
  wire [63:0] _T_213 = _T_212 | _T_208; // @[Mux.scala 27:72]
  wire [63:0] _T_214 = _T_213 | _T_30; // @[Mux.scala 27:72]
  wire  _T_219 = mipcen & _T_39; // @[CSR.scala 184:42]
  wire  _T_221 = 12'h341 == io_imme; // @[Mux.scala 80:60]
  wire [63:0] _T_222 = _T_221 ? mepcins : 64'h0; // @[Mux.scala 80:57]
  wire  _T_223 = 12'h342 == io_imme; // @[Mux.scala 80:60]
  wire [63:0] _T_224 = _T_223 ? mcauseins : _T_222; // @[Mux.scala 80:57]
  wire  _T_225 = 12'h305 == io_imme; // @[Mux.scala 80:60]
  wire [63:0] _T_226 = _T_225 ? mtvecins : _T_224; // @[Mux.scala 80:57]
  wire  _T_227 = 12'h300 == io_imme; // @[Mux.scala 80:60]
  wire [63:0] _T_228 = _T_227 ? mstatusins : _T_226; // @[Mux.scala 80:57]
  wire  _T_229 = 12'h304 == io_imme; // @[Mux.scala 80:60]
  wire [63:0] _T_230 = _T_229 ? mieins : _T_228; // @[Mux.scala 80:57]
  wire  _T_231 = 12'h344 == io_imme; // @[Mux.scala 80:60]
  wire  _T_235 = mieins[7] & mstatusins[3]; // @[CSR.scala 242:29]
  wire  startTimeCnt = _T_235; // @[CSR.scala 241:26 CSR.scala 242:16]
  assign io_rd = _T_231 ? mipins : _T_230; // @[CSR.scala 222:9]
  assign io_mtvec = mtvecins; // @[CSR.scala 238:12]
  assign io_mepc = mepcins; // @[CSR.scala 239:11]
  assign startTimeCnt_0 = startTimeCnt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mepcins = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mcauseins = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mtvecins = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mstatusins = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mieins = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mipins = _RAND_5[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      mepcins <= 64'h0;
    end else if (_T_40) begin
      if (_T_12) begin
        mepcins <= io_pc;
      end else begin
        mepcins <= _T_35;
      end
    end
    if (reset) begin
      mcauseins <= 64'h0;
    end else if (_T_73) begin
      if (intr) begin
        mcauseins <= 64'h8000000000000007;
      end else if (io_ecall) begin
        mcauseins <= 64'hb;
      end else begin
        mcauseins <= _T_67;
      end
    end
    if (reset) begin
      mtvecins <= 64'h0;
    end else if (_T_103) begin
      mtvecins <= mtvecval;
    end
    if (reset) begin
      mstatusins <= 64'ha00001800;
    end else if (_T_154) begin
      if (_T_12) begin
        mstatusins <= _T_117;
      end else if (io_mret) begin
        mstatusins <= _T_125;
      end else begin
        mstatusins <= _T_148;
      end
    end
    if (reset) begin
      mieins <= 64'h0;
    end else if (_T_184) begin
      mieins <= mieval;
    end
    if (reset) begin
      mipins <= 64'h0;
    end else if (_T_219) begin
      if (intr) begin
        mipins <= _T_191;
      end else begin
        mipins <= _T_214;
      end
    end
  end
endmodule
module dnpcGen(
  input         io_npcSrc,
  input  [31:0] io_pc,
  input  [31:0] io_imme,
  input  [31:0] io_rd,
  output [31:0] io_dnpc
);
  wire  _T = ~io_npcSrc; // @[dnpcGen.scala 15:28]
  wire [31:0] src1 = _T ? io_rd : io_pc; // @[dnpcGen.scala 15:17]
  assign io_dnpc = io_imme + src1; // @[dnpcGen.scala 16:11]
endmodule
module memData(
  input  [63:0] io_rdata,
  output [63:0] io_rdata_ext,
  input  [2:0]  io_memReadNum
);
  wire [55:0] _T_3 = io_rdata[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_4 = {_T_3,io_rdata[7:0]}; // @[Cat.scala 29:58]
  wire [47:0] _T_8 = io_rdata[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_9 = {_T_8,io_rdata[15:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_13 = io_rdata[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_14 = {_T_13,io_rdata[31:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_16 = {56'h0,io_rdata[7:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_18 = {48'h0,io_rdata[15:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_20 = {32'h0,io_rdata[31:0]}; // @[Cat.scala 29:58]
  wire  _T_21 = 3'h0 == io_memReadNum; // @[Mux.scala 80:60]
  wire [63:0] _T_22 = _T_21 ? _T_4 : 64'h0; // @[Mux.scala 80:57]
  wire  _T_23 = 3'h1 == io_memReadNum; // @[Mux.scala 80:60]
  wire [63:0] _T_24 = _T_23 ? _T_9 : _T_22; // @[Mux.scala 80:57]
  wire  _T_25 = 3'h2 == io_memReadNum; // @[Mux.scala 80:60]
  wire [63:0] _T_26 = _T_25 ? _T_14 : _T_24; // @[Mux.scala 80:57]
  wire  _T_27 = 3'h3 == io_memReadNum; // @[Mux.scala 80:60]
  wire [63:0] _T_28 = _T_27 ? io_rdata : _T_26; // @[Mux.scala 80:57]
  wire  _T_29 = 3'h4 == io_memReadNum; // @[Mux.scala 80:60]
  wire [63:0] _T_30 = _T_29 ? _T_16 : _T_28; // @[Mux.scala 80:57]
  wire  _T_31 = 3'h5 == io_memReadNum; // @[Mux.scala 80:60]
  wire [63:0] _T_32 = _T_31 ? _T_18 : _T_30; // @[Mux.scala 80:57]
  wire  _T_33 = 3'h6 == io_memReadNum; // @[Mux.scala 80:60]
  assign io_rdata_ext = _T_33 ? _T_20 : _T_32; // @[memData.scala 14:16]
endmodule
module execute(
  input          clock,
  input          reset,
  input  [1:0]   io_AluSrc1,
  input  [1:0]   io_AluSrc2,
  input  [4:0]   io_ALUCtrl,
  input          io_dnpcSrc,
  input  [1:0]   io_ResultSrc,
  input  [2:0]   io_memReadNum,
  input  [63:0]  io_dataId_imme,
  input  [63:0]  io_dataId_dOut1,
  input  [63:0]  io_dataId_dOut2,
  output [63:0]  io_dataId_dIn,
  input  [63:0]  io_dataId_rdDout,
  output [63:0]  io_dataOut_ALUResOut,
  output [63:0]  io_dataOut_wdata,
  input  [63:0]  io_dataOut_rdata,
  output         io_brTake,
  input  [31:0]  io_pc,
  input  [31:0]  io_snpc,
  output [31:0]  io_dnpc,
  input          io_CSRCtrlIf_csrrwen,
  input          io_CSRCtrlIf_csrswen,
  input          io_CSRCtrlIf_csrrsien,
  input          io_CSRCtrlIf_csrrcien,
  input          io_CSRCtrlIf_csrrcen,
  input          io_CSRCtrlIf_csrrwien,
  input          io_CSRCtrlIf_ecall,
  input          io_CSRCtrlIf_rfen,
  input          io_CSRCtrlIf_mepc2pc,
  input  [4:0]   io_uimm,
  input  [63:0]  io_aluResIn,
  input  [1:0]   io_forwardA,
  input  [1:0]   io_forwardB,
  input  [1:0]   io_forwardC,
  input  [63:0]  io_aluRes1,
  input  [63:0]  io_aluRes3,
  input          intrTimeCnt_0,
  output         startTimeCnt,
  output [191:0] dmaCtrl_0,
  input          blockDMA,
  input          block23,
  output         block1
);
  wire  ALU_clock; // @[execute.scala 99:19]
  wire  ALU_reset; // @[execute.scala 99:19]
  wire [63:0] ALU_io_srcA; // @[execute.scala 99:19]
  wire [63:0] ALU_io_srcB; // @[execute.scala 99:19]
  wire [4:0] ALU_io_ALUCtrl; // @[execute.scala 99:19]
  wire [63:0] ALU_io_ALUResult; // @[execute.scala 99:19]
  wire  ALU_block23_0; // @[execute.scala 99:19]
  wire  ALU_block1_0; // @[execute.scala 99:19]
  wire  csr_ins_clock; // @[execute.scala 106:23]
  wire  csr_ins_reset; // @[execute.scala 106:23]
  wire  csr_ins_io_csrrwen; // @[execute.scala 106:23]
  wire  csr_ins_io_csrswen; // @[execute.scala 106:23]
  wire  csr_ins_io_csrrsien; // @[execute.scala 106:23]
  wire  csr_ins_io_csrrcien; // @[execute.scala 106:23]
  wire  csr_ins_io_csrrcen; // @[execute.scala 106:23]
  wire  csr_ins_io_csrrwien; // @[execute.scala 106:23]
  wire  csr_ins_io_ecall; // @[execute.scala 106:23]
  wire [63:0] csr_ins_io_rs1; // @[execute.scala 106:23]
  wire [11:0] csr_ins_io_imme; // @[execute.scala 106:23]
  wire [63:0] csr_ins_io_pc; // @[execute.scala 106:23]
  wire [4:0] csr_ins_io_uimm; // @[execute.scala 106:23]
  wire [63:0] csr_ins_io_rd; // @[execute.scala 106:23]
  wire [63:0] csr_ins_io_mtvec; // @[execute.scala 106:23]
  wire [63:0] csr_ins_io_mepc; // @[execute.scala 106:23]
  wire  csr_ins_io_mret; // @[execute.scala 106:23]
  wire  csr_ins_intrTimeCnt_0; // @[execute.scala 106:23]
  wire  csr_ins_startTimeCnt_0; // @[execute.scala 106:23]
  wire  csr_ins_blockDMA_0; // @[execute.scala 106:23]
  wire  csr_ins_block23_0; // @[execute.scala 106:23]
  wire  csr_ins_block1_0; // @[execute.scala 106:23]
  wire  dnpcGenIns_io_npcSrc; // @[execute.scala 126:26]
  wire [31:0] dnpcGenIns_io_pc; // @[execute.scala 126:26]
  wire [31:0] dnpcGenIns_io_imme; // @[execute.scala 126:26]
  wire [31:0] dnpcGenIns_io_rd; // @[execute.scala 126:26]
  wire [31:0] dnpcGenIns_io_dnpc; // @[execute.scala 126:26]
  wire [63:0] memData_ins_io_rdata; // @[execute.scala 151:27]
  wire [63:0] memData_ins_io_rdata_ext; // @[execute.scala 151:27]
  wire [2:0] memData_ins_io_memReadNum; // @[execute.scala 151:27]
  wire  _T = 2'h2 == io_forwardA; // @[Mux.scala 80:60]
  wire [63:0] _T_1 = _T ? io_aluRes1 : io_dataId_dOut1; // @[Mux.scala 80:57]
  wire  _T_2 = 2'h1 == io_forwardA; // @[Mux.scala 80:60]
  wire  _T_30 = 2'h2 == io_ResultSrc; // @[Mux.scala 80:60]
  wire  _T_28 = 2'h1 == io_ResultSrc; // @[Mux.scala 80:60]
  wire [63:0] _T_29 = _T_28 ? {{32'd0}, io_snpc} : io_aluResIn; // @[Mux.scala 80:57]
  wire [63:0] dinMux = _T_30 ? memData_ins_io_rdata_ext : _T_29; // @[Mux.scala 80:57]
  wire [63:0] _T_3 = _T_2 ? dinMux : _T_1; // @[Mux.scala 80:57]
  wire  _T_4 = 2'h3 == io_forwardA; // @[Mux.scala 80:60]
  wire [63:0] dOut1 = _T_4 ? io_aluRes3 : _T_3; // @[Mux.scala 80:57]
  wire  _T_5 = 2'h0 == io_AluSrc1; // @[Mux.scala 80:60]
  wire [63:0] _T_6 = _T_5 ? dOut1 : 64'h0; // @[Mux.scala 80:57]
  wire  _T_7 = 2'h1 == io_AluSrc1; // @[Mux.scala 80:60]
  wire [63:0] _T_8 = _T_7 ? io_dataId_imme : _T_6; // @[Mux.scala 80:57]
  wire  _T_9 = 2'h2 == io_AluSrc1; // @[Mux.scala 80:60]
  wire  _T_10 = 2'h2 == io_forwardB; // @[Mux.scala 80:60]
  wire [63:0] _T_11 = _T_10 ? io_aluRes1 : io_dataId_dOut2; // @[Mux.scala 80:57]
  wire  _T_12 = 2'h1 == io_forwardB; // @[Mux.scala 80:60]
  wire [63:0] _T_13 = _T_12 ? dinMux : _T_11; // @[Mux.scala 80:57]
  wire  _T_14 = 2'h3 == io_forwardB; // @[Mux.scala 80:60]
  wire [63:0] dOut2 = _T_14 ? io_aluRes3 : _T_13; // @[Mux.scala 80:57]
  wire  _T_15 = 2'h0 == io_AluSrc2; // @[Mux.scala 80:60]
  wire [63:0] _T_16 = _T_15 ? dOut2 : 64'h0; // @[Mux.scala 80:57]
  wire  _T_17 = 2'h1 == io_AluSrc2; // @[Mux.scala 80:60]
  wire [63:0] _T_18 = _T_17 ? io_dataId_imme : _T_16; // @[Mux.scala 80:57]
  wire  _T_19 = 2'h2 == io_AluSrc2; // @[Mux.scala 80:60]
  wire  _T_21 = io_CSRCtrlIf_ecall | intrTimeCnt_0; // @[execute.scala 137:37]
  wire [63:0] _T_22 = io_CSRCtrlIf_mepc2pc ? csr_ins_io_mepc : {{32'd0}, dnpcGenIns_io_dnpc}; // @[execute.scala 137:72]
  wire [63:0] _T_23 = _T_21 ? csr_ins_io_mtvec : _T_22; // @[execute.scala 137:17]
  wire  _T_31 = 2'h2 == io_forwardC; // @[Mux.scala 80:60]
  wire [63:0] _T_32 = _T_31 ? io_aluRes1 : io_dataId_rdDout; // @[Mux.scala 80:57]
  wire  _T_33 = 2'h1 == io_forwardC; // @[Mux.scala 80:60]
  wire [63:0] _T_34 = _T_33 ? dinMux : _T_32; // @[Mux.scala 80:57]
  wire  _T_35 = 2'h3 == io_forwardC; // @[Mux.scala 80:60]
  wire [63:0] dmaLen = _T_35 ? io_aluRes3 : _T_34; // @[Mux.scala 80:57]
  wire [191:0] _T_37 = {dmaLen,dOut2,dOut1}; // @[Cat.scala 29:58]
  wire [191:0] dmaCtrl = _T_37; // @[execute.scala 183:21 execute.scala 184:11]
  ALU ALU ( // @[execute.scala 99:19]
    .clock(ALU_clock),
    .reset(ALU_reset),
    .io_srcA(ALU_io_srcA),
    .io_srcB(ALU_io_srcB),
    .io_ALUCtrl(ALU_io_ALUCtrl),
    .io_ALUResult(ALU_io_ALUResult),
    .block23_0(ALU_block23_0),
    .block1_0(ALU_block1_0)
  );
  CSR csr_ins ( // @[execute.scala 106:23]
    .clock(csr_ins_clock),
    .reset(csr_ins_reset),
    .io_csrrwen(csr_ins_io_csrrwen),
    .io_csrswen(csr_ins_io_csrswen),
    .io_csrrsien(csr_ins_io_csrrsien),
    .io_csrrcien(csr_ins_io_csrrcien),
    .io_csrrcen(csr_ins_io_csrrcen),
    .io_csrrwien(csr_ins_io_csrrwien),
    .io_ecall(csr_ins_io_ecall),
    .io_rs1(csr_ins_io_rs1),
    .io_imme(csr_ins_io_imme),
    .io_pc(csr_ins_io_pc),
    .io_uimm(csr_ins_io_uimm),
    .io_rd(csr_ins_io_rd),
    .io_mtvec(csr_ins_io_mtvec),
    .io_mepc(csr_ins_io_mepc),
    .io_mret(csr_ins_io_mret),
    .intrTimeCnt_0(csr_ins_intrTimeCnt_0),
    .startTimeCnt_0(csr_ins_startTimeCnt_0),
    .blockDMA_0(csr_ins_blockDMA_0),
    .block23_0(csr_ins_block23_0),
    .block1_0(csr_ins_block1_0)
  );
  dnpcGen dnpcGenIns ( // @[execute.scala 126:26]
    .io_npcSrc(dnpcGenIns_io_npcSrc),
    .io_pc(dnpcGenIns_io_pc),
    .io_imme(dnpcGenIns_io_imme),
    .io_rd(dnpcGenIns_io_rd),
    .io_dnpc(dnpcGenIns_io_dnpc)
  );
  memData memData_ins ( // @[execute.scala 151:27]
    .io_rdata(memData_ins_io_rdata),
    .io_rdata_ext(memData_ins_io_rdata_ext),
    .io_memReadNum(memData_ins_io_memReadNum)
  );
  assign io_dataId_dIn = _T_30 ? memData_ins_io_rdata_ext : _T_29; // @[execute.scala 168:17]
  assign io_dataOut_ALUResOut = io_CSRCtrlIf_rfen ? csr_ins_io_rd : ALU_io_ALUResult; // @[execute.scala 123:24]
  assign io_dataOut_wdata = _T_14 ? io_aluRes3 : _T_13; // @[execute.scala 124:20]
  assign io_brTake = ALU_io_ALUResult[0]; // @[execute.scala 139:13]
  assign io_dnpc = _T_23[31:0]; // @[execute.scala 137:11]
  assign startTimeCnt = csr_ins_startTimeCnt_0;
  assign dmaCtrl_0 = dmaCtrl;
  assign block1 = ALU_block1_0;
  assign ALU_clock = clock;
  assign ALU_reset = reset;
  assign ALU_io_srcA = _T_9 ? {{32'd0}, io_pc} : _T_8; // @[execute.scala 100:15]
  assign ALU_io_srcB = _T_19 ? {{32'd0}, io_pc} : _T_18; // @[execute.scala 101:15]
  assign ALU_io_ALUCtrl = io_ALUCtrl; // @[execute.scala 102:18]
  assign ALU_block23_0 = block23;
  assign csr_ins_clock = clock;
  assign csr_ins_reset = reset;
  assign csr_ins_io_csrrwen = io_CSRCtrlIf_csrrwen; // @[execute.scala 107:22]
  assign csr_ins_io_csrswen = io_CSRCtrlIf_csrswen; // @[execute.scala 108:22]
  assign csr_ins_io_csrrsien = io_CSRCtrlIf_csrrsien; // @[execute.scala 109:23]
  assign csr_ins_io_csrrcien = io_CSRCtrlIf_csrrcien; // @[execute.scala 110:23]
  assign csr_ins_io_csrrcen = io_CSRCtrlIf_csrrcen; // @[execute.scala 111:22]
  assign csr_ins_io_csrrwien = io_CSRCtrlIf_csrrwien; // @[execute.scala 112:23]
  assign csr_ins_io_ecall = io_CSRCtrlIf_ecall; // @[execute.scala 113:20]
  assign csr_ins_io_rs1 = _T_4 ? io_aluRes3 : _T_3; // @[execute.scala 115:18]
  assign csr_ins_io_imme = io_dataId_imme[11:0]; // @[execute.scala 116:19]
  assign csr_ins_io_pc = {{32'd0}, io_pc}; // @[execute.scala 117:17]
  assign csr_ins_io_uimm = io_uimm; // @[execute.scala 118:19]
  assign csr_ins_io_mret = io_CSRCtrlIf_mepc2pc; // @[execute.scala 119:19]
  assign csr_ins_intrTimeCnt_0 = intrTimeCnt_0;
  assign csr_ins_blockDMA_0 = blockDMA;
  assign csr_ins_block23_0 = block23;
  assign csr_ins_block1_0 = block1;
  assign dnpcGenIns_io_npcSrc = io_dnpcSrc; // @[execute.scala 131:24]
  assign dnpcGenIns_io_pc = io_pc; // @[execute.scala 127:20]
  assign dnpcGenIns_io_imme = io_dataId_imme[31:0]; // @[execute.scala 128:22]
  assign dnpcGenIns_io_rd = dOut1[31:0]; // @[execute.scala 130:20]
  assign memData_ins_io_rdata = io_dataOut_rdata; // @[execute.scala 153:24]
  assign memData_ins_io_memReadNum = io_memReadNum; // @[execute.scala 152:29]
endmodule
module hazard(
  input        io_regEnEXMEM,
  input  [4:0] io_rdEXMEM,
  input  [4:0] io_rs1IDEX,
  input  [4:0] io_rs2IDEX,
  input        io_regEnMEMWB,
  input  [4:0] io_rdMEMWB,
  input        io_regEnWBEND,
  input  [4:0] io_rdWBEND,
  output [1:0] io_forwardA,
  output [1:0] io_forwardB,
  output [1:0] io_forwardC,
  input  [4:0] io_rs1IFID,
  input  [4:0] io_rs2IFID,
  input  [4:0] io_rdIDEX,
  input  [1:0] io_resSrc,
  output       io_loadHazard
);
  wire  _T = io_rdEXMEM == io_rs1IDEX; // @[hazard.scala 39:48]
  wire  _T_1 = io_regEnEXMEM & _T; // @[hazard.scala 39:35]
  wire  _T_2 = io_rs1IDEX != 5'h0; // @[hazard.scala 39:76]
  wire  forwardAOne = _T_1 & _T_2; // @[hazard.scala 39:63]
  wire  _T_3 = io_rdMEMWB == io_rs1IDEX; // @[hazard.scala 40:49]
  wire  _T_4 = io_regEnMEMWB & _T_3; // @[hazard.scala 40:35]
  wire  _T_6 = _T_4 & _T_2; // @[hazard.scala 40:64]
  wire  _T_7 = io_rdEXMEM != io_rs1IDEX; // @[hazard.scala 40:97]
  wire  _T_8 = ~io_regEnEXMEM; // @[hazard.scala 40:115]
  wire  _T_9 = _T_7 | _T_8; // @[hazard.scala 40:112]
  wire  forwardATwo = _T_6 & _T_9; // @[hazard.scala 40:84]
  wire  _T_10 = io_rdWBEND == io_rs1IDEX; // @[hazard.scala 41:51]
  wire  _T_11 = io_regEnWBEND & _T_10; // @[hazard.scala 41:37]
  wire  forwardAThree = _T_11 & _T_2; // @[hazard.scala 41:66]
  wire [1:0] _T_13 = forwardAThree ? 2'h3 : 2'h0; // @[hazard.scala 42:75]
  wire [1:0] _T_14 = forwardATwo ? 2'h1 : _T_13; // @[hazard.scala 42:47]
  wire  _T_16 = io_rdEXMEM == io_rs2IDEX; // @[hazard.scala 44:48]
  wire  _T_17 = io_regEnEXMEM & _T_16; // @[hazard.scala 44:35]
  wire  _T_18 = io_rs2IDEX != 5'h0; // @[hazard.scala 44:76]
  wire  forwardBOne = _T_17 & _T_18; // @[hazard.scala 44:63]
  wire  _T_19 = io_rdMEMWB == io_rs2IDEX; // @[hazard.scala 45:49]
  wire  _T_20 = io_regEnMEMWB & _T_19; // @[hazard.scala 45:35]
  wire  _T_22 = _T_20 & _T_18; // @[hazard.scala 45:64]
  wire  _T_23 = io_rdEXMEM != io_rs2IDEX; // @[hazard.scala 45:97]
  wire  _T_25 = _T_23 | _T_8; // @[hazard.scala 45:112]
  wire  forwardBTwo = _T_22 & _T_25; // @[hazard.scala 45:84]
  wire  _T_26 = io_rdWBEND == io_rs2IDEX; // @[hazard.scala 46:52]
  wire  _T_27 = io_regEnWBEND & _T_26; // @[hazard.scala 46:38]
  wire  forwardBThree = _T_27 & _T_18; // @[hazard.scala 46:67]
  wire [1:0] _T_29 = forwardBThree ? 2'h3 : 2'h0; // @[hazard.scala 47:75]
  wire [1:0] _T_30 = forwardBTwo ? 2'h1 : _T_29; // @[hazard.scala 47:47]
  wire  _T_32 = io_rdEXMEM == io_rdIDEX; // @[hazard.scala 50:49]
  wire  _T_33 = io_regEnEXMEM & _T_32; // @[hazard.scala 50:35]
  wire  _T_34 = io_rdIDEX != 5'h0; // @[hazard.scala 50:76]
  wire  forwardCOne = _T_33 & _T_34; // @[hazard.scala 50:63]
  wire  _T_35 = io_rdMEMWB == io_rdIDEX; // @[hazard.scala 51:49]
  wire  _T_36 = io_regEnMEMWB & _T_35; // @[hazard.scala 51:35]
  wire  _T_38 = _T_36 & _T_34; // @[hazard.scala 51:63]
  wire  _T_39 = io_rdEXMEM != io_rdIDEX; // @[hazard.scala 51:99]
  wire  _T_41 = _T_39 | _T_8; // @[hazard.scala 51:113]
  wire  forwardCTwo = _T_38 & _T_41; // @[hazard.scala 51:84]
  wire  _T_42 = io_rdWBEND == io_rdIDEX; // @[hazard.scala 52:51]
  wire  _T_43 = io_regEnWBEND & _T_42; // @[hazard.scala 52:37]
  wire  forwardCThree = _T_43 & _T_34; // @[hazard.scala 52:65]
  wire [1:0] _T_45 = forwardCThree ? 2'h3 : 2'h0; // @[hazard.scala 53:75]
  wire [1:0] _T_46 = forwardCTwo ? 2'h1 : _T_45; // @[hazard.scala 53:48]
  wire  _T_48 = io_rs1IFID == io_rdIDEX; // @[hazard.scala 58:32]
  wire  _T_49 = io_rs2IFID == io_rdIDEX; // @[hazard.scala 58:59]
  wire  _T_50 = _T_48 | _T_49; // @[hazard.scala 58:46]
  wire  _T_51 = io_resSrc == 2'h2; // @[hazard.scala 58:87]
  assign io_forwardA = forwardAOne ? 2'h2 : _T_14; // @[hazard.scala 42:15]
  assign io_forwardB = forwardBOne ? 2'h2 : _T_30; // @[hazard.scala 47:15]
  assign io_forwardC = forwardCOne ? 2'h2 : _T_46; // @[hazard.scala 53:15]
  assign io_loadHazard = _T_50 & _T_51; // @[hazard.scala 58:17]
endmodule
module preCell(
  input         clock,
  input         reset,
  input         io_cen,
  input         io_jump,
  input  [31:0] io_dnpcIn,
  output [31:0] io_dnpcOut,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _T = io_cen & io_jump; // @[preCell.scala 17:48]
  reg [31:0] dnpcReg; // @[Reg.scala 27:20]
  wire  takenV = dnpcReg == io_dnpcIn; // @[preCell.scala 22:24]
  reg [1:0] stateWire; // @[Reg.scala 27:20]
  wire  _T_1 = 2'h1 == stateWire; // @[Mux.scala 80:60]
  wire  _T_3 = 2'h2 == stateWire; // @[Mux.scala 80:60]
  wire  _T_5 = 2'h3 == stateWire; // @[Mux.scala 80:60]
  wire  _T_8 = stateWire == 2'h2; // @[preCell.scala 44:25]
  wire  _T_9 = stateWire == 2'h3; // @[preCell.scala 44:49]
  assign io_dnpcOut = dnpcReg; // @[preCell.scala 43:14]
  assign io_valid = _T_8 | _T_9; // @[preCell.scala 44:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dnpcReg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  stateWire = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      dnpcReg <= 32'h0;
    end else if (_T) begin
      dnpcReg <= io_dnpcIn;
    end
    if (reset) begin
      stateWire <= 2'h0;
    end else if (io_cen) begin
      if (_T_5) begin
        if (takenV) begin
          stateWire <= 2'h3;
        end else begin
          stateWire <= 2'h2;
        end
      end else if (_T_3) begin
        if (takenV) begin
          stateWire <= 2'h3;
        end else begin
          stateWire <= 2'h1;
        end
      end else if (_T_1) begin
        if (takenV) begin
          stateWire <= 2'h2;
        end else begin
          stateWire <= 2'h0;
        end
      end else if (takenV) begin
        stateWire <= 2'h1;
      end else begin
        stateWire <= 2'h0;
      end
    end
  end
endmodule
module preBranch(
  input         clock,
  input         reset,
  input         io_exjump,
  input  [31:0] io_ifpc,
  input  [31:0] io_expc,
  input  [31:0] io_exdpc,
  output [31:0] io_ifdnpc,
  output        io_ifjump,
  input         block23_0,
  input         block1_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  wire  precelList_0_clock; // @[preBranch.scala 30:45]
  wire  precelList_0_reset; // @[preBranch.scala 30:45]
  wire  precelList_0_io_cen; // @[preBranch.scala 30:45]
  wire  precelList_0_io_jump; // @[preBranch.scala 30:45]
  wire [31:0] precelList_0_io_dnpcIn; // @[preBranch.scala 30:45]
  wire [31:0] precelList_0_io_dnpcOut; // @[preBranch.scala 30:45]
  wire  precelList_0_io_valid; // @[preBranch.scala 30:45]
  wire  precelList_1_clock; // @[preBranch.scala 30:45]
  wire  precelList_1_reset; // @[preBranch.scala 30:45]
  wire  precelList_1_io_cen; // @[preBranch.scala 30:45]
  wire  precelList_1_io_jump; // @[preBranch.scala 30:45]
  wire [31:0] precelList_1_io_dnpcIn; // @[preBranch.scala 30:45]
  wire [31:0] precelList_1_io_dnpcOut; // @[preBranch.scala 30:45]
  wire  precelList_1_io_valid; // @[preBranch.scala 30:45]
  wire  precelList_2_clock; // @[preBranch.scala 30:45]
  wire  precelList_2_reset; // @[preBranch.scala 30:45]
  wire  precelList_2_io_cen; // @[preBranch.scala 30:45]
  wire  precelList_2_io_jump; // @[preBranch.scala 30:45]
  wire [31:0] precelList_2_io_dnpcIn; // @[preBranch.scala 30:45]
  wire [31:0] precelList_2_io_dnpcOut; // @[preBranch.scala 30:45]
  wire  precelList_2_io_valid; // @[preBranch.scala 30:45]
  wire  precelList_3_clock; // @[preBranch.scala 30:45]
  wire  precelList_3_reset; // @[preBranch.scala 30:45]
  wire  precelList_3_io_cen; // @[preBranch.scala 30:45]
  wire  precelList_3_io_jump; // @[preBranch.scala 30:45]
  wire [31:0] precelList_3_io_dnpcIn; // @[preBranch.scala 30:45]
  wire [31:0] precelList_3_io_dnpcOut; // @[preBranch.scala 30:45]
  wire  precelList_3_io_valid; // @[preBranch.scala 30:45]
  wire  precelList_4_clock; // @[preBranch.scala 30:45]
  wire  precelList_4_reset; // @[preBranch.scala 30:45]
  wire  precelList_4_io_cen; // @[preBranch.scala 30:45]
  wire  precelList_4_io_jump; // @[preBranch.scala 30:45]
  wire [31:0] precelList_4_io_dnpcIn; // @[preBranch.scala 30:45]
  wire [31:0] precelList_4_io_dnpcOut; // @[preBranch.scala 30:45]
  wire  precelList_4_io_valid; // @[preBranch.scala 30:45]
  wire  precelList_5_clock; // @[preBranch.scala 30:45]
  wire  precelList_5_reset; // @[preBranch.scala 30:45]
  wire  precelList_5_io_cen; // @[preBranch.scala 30:45]
  wire  precelList_5_io_jump; // @[preBranch.scala 30:45]
  wire [31:0] precelList_5_io_dnpcIn; // @[preBranch.scala 30:45]
  wire [31:0] precelList_5_io_dnpcOut; // @[preBranch.scala 30:45]
  wire  precelList_5_io_valid; // @[preBranch.scala 30:45]
  wire  precelList_6_clock; // @[preBranch.scala 30:45]
  wire  precelList_6_reset; // @[preBranch.scala 30:45]
  wire  precelList_6_io_cen; // @[preBranch.scala 30:45]
  wire  precelList_6_io_jump; // @[preBranch.scala 30:45]
  wire [31:0] precelList_6_io_dnpcIn; // @[preBranch.scala 30:45]
  wire [31:0] precelList_6_io_dnpcOut; // @[preBranch.scala 30:45]
  wire  precelList_6_io_valid; // @[preBranch.scala 30:45]
  wire  precelList_7_clock; // @[preBranch.scala 30:45]
  wire  precelList_7_reset; // @[preBranch.scala 30:45]
  wire  precelList_7_io_cen; // @[preBranch.scala 30:45]
  wire  precelList_7_io_jump; // @[preBranch.scala 30:45]
  wire [31:0] precelList_7_io_dnpcIn; // @[preBranch.scala 30:45]
  wire [31:0] precelList_7_io_dnpcOut; // @[preBranch.scala 30:45]
  wire  precelList_7_io_valid; // @[preBranch.scala 30:45]
  wire  precelList_8_clock; // @[preBranch.scala 30:45]
  wire  precelList_8_reset; // @[preBranch.scala 30:45]
  wire  precelList_8_io_cen; // @[preBranch.scala 30:45]
  wire  precelList_8_io_jump; // @[preBranch.scala 30:45]
  wire [31:0] precelList_8_io_dnpcIn; // @[preBranch.scala 30:45]
  wire [31:0] precelList_8_io_dnpcOut; // @[preBranch.scala 30:45]
  wire  precelList_8_io_valid; // @[preBranch.scala 30:45]
  wire  precelList_9_clock; // @[preBranch.scala 30:45]
  wire  precelList_9_reset; // @[preBranch.scala 30:45]
  wire  precelList_9_io_cen; // @[preBranch.scala 30:45]
  wire  precelList_9_io_jump; // @[preBranch.scala 30:45]
  wire [31:0] precelList_9_io_dnpcIn; // @[preBranch.scala 30:45]
  wire [31:0] precelList_9_io_dnpcOut; // @[preBranch.scala 30:45]
  wire  precelList_9_io_valid; // @[preBranch.scala 30:45]
  wire  precelList_10_clock; // @[preBranch.scala 30:45]
  wire  precelList_10_reset; // @[preBranch.scala 30:45]
  wire  precelList_10_io_cen; // @[preBranch.scala 30:45]
  wire  precelList_10_io_jump; // @[preBranch.scala 30:45]
  wire [31:0] precelList_10_io_dnpcIn; // @[preBranch.scala 30:45]
  wire [31:0] precelList_10_io_dnpcOut; // @[preBranch.scala 30:45]
  wire  precelList_10_io_valid; // @[preBranch.scala 30:45]
  wire  precelList_11_clock; // @[preBranch.scala 30:45]
  wire  precelList_11_reset; // @[preBranch.scala 30:45]
  wire  precelList_11_io_cen; // @[preBranch.scala 30:45]
  wire  precelList_11_io_jump; // @[preBranch.scala 30:45]
  wire [31:0] precelList_11_io_dnpcIn; // @[preBranch.scala 30:45]
  wire [31:0] precelList_11_io_dnpcOut; // @[preBranch.scala 30:45]
  wire  precelList_11_io_valid; // @[preBranch.scala 30:45]
  wire  precelList_12_clock; // @[preBranch.scala 30:45]
  wire  precelList_12_reset; // @[preBranch.scala 30:45]
  wire  precelList_12_io_cen; // @[preBranch.scala 30:45]
  wire  precelList_12_io_jump; // @[preBranch.scala 30:45]
  wire [31:0] precelList_12_io_dnpcIn; // @[preBranch.scala 30:45]
  wire [31:0] precelList_12_io_dnpcOut; // @[preBranch.scala 30:45]
  wire  precelList_12_io_valid; // @[preBranch.scala 30:45]
  wire  precelList_13_clock; // @[preBranch.scala 30:45]
  wire  precelList_13_reset; // @[preBranch.scala 30:45]
  wire  precelList_13_io_cen; // @[preBranch.scala 30:45]
  wire  precelList_13_io_jump; // @[preBranch.scala 30:45]
  wire [31:0] precelList_13_io_dnpcIn; // @[preBranch.scala 30:45]
  wire [31:0] precelList_13_io_dnpcOut; // @[preBranch.scala 30:45]
  wire  precelList_13_io_valid; // @[preBranch.scala 30:45]
  wire  precelList_14_clock; // @[preBranch.scala 30:45]
  wire  precelList_14_reset; // @[preBranch.scala 30:45]
  wire  precelList_14_io_cen; // @[preBranch.scala 30:45]
  wire  precelList_14_io_jump; // @[preBranch.scala 30:45]
  wire [31:0] precelList_14_io_dnpcIn; // @[preBranch.scala 30:45]
  wire [31:0] precelList_14_io_dnpcOut; // @[preBranch.scala 30:45]
  wire  precelList_14_io_valid; // @[preBranch.scala 30:45]
  wire  precelList_15_clock; // @[preBranch.scala 30:45]
  wire  precelList_15_reset; // @[preBranch.scala 30:45]
  wire  precelList_15_io_cen; // @[preBranch.scala 30:45]
  wire  precelList_15_io_jump; // @[preBranch.scala 30:45]
  wire [31:0] precelList_15_io_dnpcIn; // @[preBranch.scala 30:45]
  wire [31:0] precelList_15_io_dnpcOut; // @[preBranch.scala 30:45]
  wire  precelList_15_io_valid; // @[preBranch.scala 30:45]
  wire  block = block1_0 | block23_0; // @[preBranch.scala 27:33]
  reg [31:0] pcList_0; // @[Reg.scala 27:20]
  wire  _T_1 = io_expc == pcList_0; // @[preBranch.scala 36:27]
  reg  vList_0; // @[Reg.scala 27:20]
  wire  hitList_0 = _T_1 & vList_0; // @[preBranch.scala 36:41]
  reg [31:0] pcList_1; // @[Reg.scala 27:20]
  wire  _T_3 = io_expc == pcList_1; // @[preBranch.scala 36:27]
  reg  vList_1; // @[Reg.scala 27:20]
  wire  hitList_1 = _T_3 & vList_1; // @[preBranch.scala 36:41]
  reg [31:0] pcList_2; // @[Reg.scala 27:20]
  wire  _T_5 = io_expc == pcList_2; // @[preBranch.scala 36:27]
  reg  vList_2; // @[Reg.scala 27:20]
  wire  hitList_2 = _T_5 & vList_2; // @[preBranch.scala 36:41]
  reg [31:0] pcList_3; // @[Reg.scala 27:20]
  wire  _T_7 = io_expc == pcList_3; // @[preBranch.scala 36:27]
  reg  vList_3; // @[Reg.scala 27:20]
  wire  hitList_3 = _T_7 & vList_3; // @[preBranch.scala 36:41]
  reg [31:0] pcList_4; // @[Reg.scala 27:20]
  wire  _T_9 = io_expc == pcList_4; // @[preBranch.scala 36:27]
  reg  vList_4; // @[Reg.scala 27:20]
  wire  hitList_4 = _T_9 & vList_4; // @[preBranch.scala 36:41]
  reg [31:0] pcList_5; // @[Reg.scala 27:20]
  wire  _T_11 = io_expc == pcList_5; // @[preBranch.scala 36:27]
  reg  vList_5; // @[Reg.scala 27:20]
  wire  hitList_5 = _T_11 & vList_5; // @[preBranch.scala 36:41]
  reg [31:0] pcList_6; // @[Reg.scala 27:20]
  wire  _T_13 = io_expc == pcList_6; // @[preBranch.scala 36:27]
  reg  vList_6; // @[Reg.scala 27:20]
  wire  hitList_6 = _T_13 & vList_6; // @[preBranch.scala 36:41]
  reg [31:0] pcList_7; // @[Reg.scala 27:20]
  wire  _T_15 = io_expc == pcList_7; // @[preBranch.scala 36:27]
  reg  vList_7; // @[Reg.scala 27:20]
  wire  hitList_7 = _T_15 & vList_7; // @[preBranch.scala 36:41]
  reg [31:0] pcList_8; // @[Reg.scala 27:20]
  wire  _T_17 = io_expc == pcList_8; // @[preBranch.scala 36:27]
  reg  vList_8; // @[Reg.scala 27:20]
  wire  hitList_8 = _T_17 & vList_8; // @[preBranch.scala 36:41]
  reg [31:0] pcList_9; // @[Reg.scala 27:20]
  wire  _T_19 = io_expc == pcList_9; // @[preBranch.scala 36:27]
  reg  vList_9; // @[Reg.scala 27:20]
  wire  hitList_9 = _T_19 & vList_9; // @[preBranch.scala 36:41]
  reg [31:0] pcList_10; // @[Reg.scala 27:20]
  wire  _T_21 = io_expc == pcList_10; // @[preBranch.scala 36:27]
  reg  vList_10; // @[Reg.scala 27:20]
  wire  hitList_10 = _T_21 & vList_10; // @[preBranch.scala 36:41]
  reg [31:0] pcList_11; // @[Reg.scala 27:20]
  wire  _T_23 = io_expc == pcList_11; // @[preBranch.scala 36:27]
  reg  vList_11; // @[Reg.scala 27:20]
  wire  hitList_11 = _T_23 & vList_11; // @[preBranch.scala 36:41]
  reg [31:0] pcList_12; // @[Reg.scala 27:20]
  wire  _T_25 = io_expc == pcList_12; // @[preBranch.scala 36:27]
  reg  vList_12; // @[Reg.scala 27:20]
  wire  hitList_12 = _T_25 & vList_12; // @[preBranch.scala 36:41]
  reg [31:0] pcList_13; // @[Reg.scala 27:20]
  wire  _T_27 = io_expc == pcList_13; // @[preBranch.scala 36:27]
  reg  vList_13; // @[Reg.scala 27:20]
  wire  hitList_13 = _T_27 & vList_13; // @[preBranch.scala 36:41]
  reg [31:0] pcList_14; // @[Reg.scala 27:20]
  wire  _T_29 = io_expc == pcList_14; // @[preBranch.scala 36:27]
  reg  vList_14; // @[Reg.scala 27:20]
  wire  hitList_14 = _T_29 & vList_14; // @[preBranch.scala 36:41]
  reg [31:0] pcList_15; // @[Reg.scala 27:20]
  wire  _T_31 = io_expc == pcList_15; // @[preBranch.scala 36:27]
  reg  vList_15; // @[Reg.scala 27:20]
  wire  hitList_15 = _T_31 & vList_15; // @[preBranch.scala 36:41]
  wire  _T_34 = hitList_0 | hitList_1; // @[preBranch.scala 38:51]
  wire  _T_35 = _T_34 | hitList_2; // @[preBranch.scala 38:51]
  wire  _T_36 = _T_35 | hitList_3; // @[preBranch.scala 38:51]
  wire  _T_37 = _T_36 | hitList_4; // @[preBranch.scala 38:51]
  wire  _T_38 = _T_37 | hitList_5; // @[preBranch.scala 38:51]
  wire  _T_39 = _T_38 | hitList_6; // @[preBranch.scala 38:51]
  wire  _T_40 = _T_39 | hitList_7; // @[preBranch.scala 38:51]
  wire  _T_41 = _T_40 | hitList_8; // @[preBranch.scala 38:51]
  wire  _T_42 = _T_41 | hitList_9; // @[preBranch.scala 38:51]
  wire  _T_43 = _T_42 | hitList_10; // @[preBranch.scala 38:51]
  wire  _T_44 = _T_43 | hitList_11; // @[preBranch.scala 38:51]
  wire  _T_45 = _T_44 | hitList_12; // @[preBranch.scala 38:51]
  wire  _T_46 = _T_45 | hitList_13; // @[preBranch.scala 38:51]
  wire  _T_47 = _T_46 | hitList_14; // @[preBranch.scala 38:51]
  wire  hit = _T_47 | hitList_15; // @[preBranch.scala 38:51]
  reg [3:0] cnt; // @[Reg.scala 27:20]
  wire [3:0] _T_49 = cnt + 4'h1; // @[preBranch.scala 41:25]
  wire  _T_50 = ~hit; // @[preBranch.scala 41:40]
  wire  _T_51 = _T_50 & io_exjump; // @[preBranch.scala 41:45]
  wire  _T_52 = ~block; // @[preBranch.scala 41:61]
  wire  _T_53 = _T_51 & _T_52; // @[preBranch.scala 41:58]
  wire  _T_55 = cnt == 4'h0; // @[preBranch.scala 47:62]
  wire  _T_56 = io_exjump & _T_55; // @[preBranch.scala 47:55]
  wire  _T_57 = hitList_0 | _T_56; // @[preBranch.scala 47:41]
  wire  _T_60 = ~hitList_0; // @[preBranch.scala 49:44]
  wire  _T_61 = _T_60 & io_exjump; // @[preBranch.scala 49:55]
  wire  _T_63 = _T_61 & _T_55; // @[preBranch.scala 49:67]
  wire  _T_65 = _T_63 & _T_52; // @[preBranch.scala 49:82]
  wire  _GEN_1 = _T_65 | vList_0; // @[Reg.scala 28:19]
  wire  _T_74 = cnt == 4'h1; // @[preBranch.scala 47:62]
  wire  _T_75 = io_exjump & _T_74; // @[preBranch.scala 47:55]
  wire  _T_76 = hitList_1 | _T_75; // @[preBranch.scala 47:41]
  wire  _T_79 = ~hitList_1; // @[preBranch.scala 49:44]
  wire  _T_80 = _T_79 & io_exjump; // @[preBranch.scala 49:55]
  wire  _T_82 = _T_80 & _T_74; // @[preBranch.scala 49:67]
  wire  _T_84 = _T_82 & _T_52; // @[preBranch.scala 49:82]
  wire  _GEN_3 = _T_84 | vList_1; // @[Reg.scala 28:19]
  wire  _T_93 = cnt == 4'h2; // @[preBranch.scala 47:62]
  wire  _T_94 = io_exjump & _T_93; // @[preBranch.scala 47:55]
  wire  _T_95 = hitList_2 | _T_94; // @[preBranch.scala 47:41]
  wire  _T_98 = ~hitList_2; // @[preBranch.scala 49:44]
  wire  _T_99 = _T_98 & io_exjump; // @[preBranch.scala 49:55]
  wire  _T_101 = _T_99 & _T_93; // @[preBranch.scala 49:67]
  wire  _T_103 = _T_101 & _T_52; // @[preBranch.scala 49:82]
  wire  _GEN_5 = _T_103 | vList_2; // @[Reg.scala 28:19]
  wire  _T_112 = cnt == 4'h3; // @[preBranch.scala 47:62]
  wire  _T_113 = io_exjump & _T_112; // @[preBranch.scala 47:55]
  wire  _T_114 = hitList_3 | _T_113; // @[preBranch.scala 47:41]
  wire  _T_117 = ~hitList_3; // @[preBranch.scala 49:44]
  wire  _T_118 = _T_117 & io_exjump; // @[preBranch.scala 49:55]
  wire  _T_120 = _T_118 & _T_112; // @[preBranch.scala 49:67]
  wire  _T_122 = _T_120 & _T_52; // @[preBranch.scala 49:82]
  wire  _GEN_7 = _T_122 | vList_3; // @[Reg.scala 28:19]
  wire  _T_131 = cnt == 4'h4; // @[preBranch.scala 47:62]
  wire  _T_132 = io_exjump & _T_131; // @[preBranch.scala 47:55]
  wire  _T_133 = hitList_4 | _T_132; // @[preBranch.scala 47:41]
  wire  _T_136 = ~hitList_4; // @[preBranch.scala 49:44]
  wire  _T_137 = _T_136 & io_exjump; // @[preBranch.scala 49:55]
  wire  _T_139 = _T_137 & _T_131; // @[preBranch.scala 49:67]
  wire  _T_141 = _T_139 & _T_52; // @[preBranch.scala 49:82]
  wire  _GEN_9 = _T_141 | vList_4; // @[Reg.scala 28:19]
  wire  _T_150 = cnt == 4'h5; // @[preBranch.scala 47:62]
  wire  _T_151 = io_exjump & _T_150; // @[preBranch.scala 47:55]
  wire  _T_152 = hitList_5 | _T_151; // @[preBranch.scala 47:41]
  wire  _T_155 = ~hitList_5; // @[preBranch.scala 49:44]
  wire  _T_156 = _T_155 & io_exjump; // @[preBranch.scala 49:55]
  wire  _T_158 = _T_156 & _T_150; // @[preBranch.scala 49:67]
  wire  _T_160 = _T_158 & _T_52; // @[preBranch.scala 49:82]
  wire  _GEN_11 = _T_160 | vList_5; // @[Reg.scala 28:19]
  wire  _T_169 = cnt == 4'h6; // @[preBranch.scala 47:62]
  wire  _T_170 = io_exjump & _T_169; // @[preBranch.scala 47:55]
  wire  _T_171 = hitList_6 | _T_170; // @[preBranch.scala 47:41]
  wire  _T_174 = ~hitList_6; // @[preBranch.scala 49:44]
  wire  _T_175 = _T_174 & io_exjump; // @[preBranch.scala 49:55]
  wire  _T_177 = _T_175 & _T_169; // @[preBranch.scala 49:67]
  wire  _T_179 = _T_177 & _T_52; // @[preBranch.scala 49:82]
  wire  _GEN_13 = _T_179 | vList_6; // @[Reg.scala 28:19]
  wire  _T_188 = cnt == 4'h7; // @[preBranch.scala 47:62]
  wire  _T_189 = io_exjump & _T_188; // @[preBranch.scala 47:55]
  wire  _T_190 = hitList_7 | _T_189; // @[preBranch.scala 47:41]
  wire  _T_193 = ~hitList_7; // @[preBranch.scala 49:44]
  wire  _T_194 = _T_193 & io_exjump; // @[preBranch.scala 49:55]
  wire  _T_196 = _T_194 & _T_188; // @[preBranch.scala 49:67]
  wire  _T_198 = _T_196 & _T_52; // @[preBranch.scala 49:82]
  wire  _GEN_15 = _T_198 | vList_7; // @[Reg.scala 28:19]
  wire  _T_207 = cnt == 4'h8; // @[preBranch.scala 47:62]
  wire  _T_208 = io_exjump & _T_207; // @[preBranch.scala 47:55]
  wire  _T_209 = hitList_8 | _T_208; // @[preBranch.scala 47:41]
  wire  _T_212 = ~hitList_8; // @[preBranch.scala 49:44]
  wire  _T_213 = _T_212 & io_exjump; // @[preBranch.scala 49:55]
  wire  _T_215 = _T_213 & _T_207; // @[preBranch.scala 49:67]
  wire  _T_217 = _T_215 & _T_52; // @[preBranch.scala 49:82]
  wire  _GEN_17 = _T_217 | vList_8; // @[Reg.scala 28:19]
  wire  _T_226 = cnt == 4'h9; // @[preBranch.scala 47:62]
  wire  _T_227 = io_exjump & _T_226; // @[preBranch.scala 47:55]
  wire  _T_228 = hitList_9 | _T_227; // @[preBranch.scala 47:41]
  wire  _T_231 = ~hitList_9; // @[preBranch.scala 49:44]
  wire  _T_232 = _T_231 & io_exjump; // @[preBranch.scala 49:55]
  wire  _T_234 = _T_232 & _T_226; // @[preBranch.scala 49:67]
  wire  _T_236 = _T_234 & _T_52; // @[preBranch.scala 49:82]
  wire  _GEN_19 = _T_236 | vList_9; // @[Reg.scala 28:19]
  wire  _T_245 = cnt == 4'ha; // @[preBranch.scala 47:62]
  wire  _T_246 = io_exjump & _T_245; // @[preBranch.scala 47:55]
  wire  _T_247 = hitList_10 | _T_246; // @[preBranch.scala 47:41]
  wire  _T_250 = ~hitList_10; // @[preBranch.scala 49:44]
  wire  _T_251 = _T_250 & io_exjump; // @[preBranch.scala 49:55]
  wire  _T_253 = _T_251 & _T_245; // @[preBranch.scala 49:67]
  wire  _T_255 = _T_253 & _T_52; // @[preBranch.scala 49:82]
  wire  _GEN_21 = _T_255 | vList_10; // @[Reg.scala 28:19]
  wire  _T_264 = cnt == 4'hb; // @[preBranch.scala 47:62]
  wire  _T_265 = io_exjump & _T_264; // @[preBranch.scala 47:55]
  wire  _T_266 = hitList_11 | _T_265; // @[preBranch.scala 47:41]
  wire  _T_269 = ~hitList_11; // @[preBranch.scala 49:44]
  wire  _T_270 = _T_269 & io_exjump; // @[preBranch.scala 49:55]
  wire  _T_272 = _T_270 & _T_264; // @[preBranch.scala 49:67]
  wire  _T_274 = _T_272 & _T_52; // @[preBranch.scala 49:82]
  wire  _GEN_23 = _T_274 | vList_11; // @[Reg.scala 28:19]
  wire  _T_283 = cnt == 4'hc; // @[preBranch.scala 47:62]
  wire  _T_284 = io_exjump & _T_283; // @[preBranch.scala 47:55]
  wire  _T_285 = hitList_12 | _T_284; // @[preBranch.scala 47:41]
  wire  _T_288 = ~hitList_12; // @[preBranch.scala 49:44]
  wire  _T_289 = _T_288 & io_exjump; // @[preBranch.scala 49:55]
  wire  _T_291 = _T_289 & _T_283; // @[preBranch.scala 49:67]
  wire  _T_293 = _T_291 & _T_52; // @[preBranch.scala 49:82]
  wire  _GEN_25 = _T_293 | vList_12; // @[Reg.scala 28:19]
  wire  _T_302 = cnt == 4'hd; // @[preBranch.scala 47:62]
  wire  _T_303 = io_exjump & _T_302; // @[preBranch.scala 47:55]
  wire  _T_304 = hitList_13 | _T_303; // @[preBranch.scala 47:41]
  wire  _T_307 = ~hitList_13; // @[preBranch.scala 49:44]
  wire  _T_308 = _T_307 & io_exjump; // @[preBranch.scala 49:55]
  wire  _T_310 = _T_308 & _T_302; // @[preBranch.scala 49:67]
  wire  _T_312 = _T_310 & _T_52; // @[preBranch.scala 49:82]
  wire  _GEN_27 = _T_312 | vList_13; // @[Reg.scala 28:19]
  wire  _T_321 = cnt == 4'he; // @[preBranch.scala 47:62]
  wire  _T_322 = io_exjump & _T_321; // @[preBranch.scala 47:55]
  wire  _T_323 = hitList_14 | _T_322; // @[preBranch.scala 47:41]
  wire  _T_326 = ~hitList_14; // @[preBranch.scala 49:44]
  wire  _T_327 = _T_326 & io_exjump; // @[preBranch.scala 49:55]
  wire  _T_329 = _T_327 & _T_321; // @[preBranch.scala 49:67]
  wire  _T_331 = _T_329 & _T_52; // @[preBranch.scala 49:82]
  wire  _GEN_29 = _T_331 | vList_14; // @[Reg.scala 28:19]
  wire  _T_340 = cnt == 4'hf; // @[preBranch.scala 47:62]
  wire  _T_341 = io_exjump & _T_340; // @[preBranch.scala 47:55]
  wire  _T_342 = hitList_15 | _T_341; // @[preBranch.scala 47:41]
  wire  _T_345 = ~hitList_15; // @[preBranch.scala 49:44]
  wire  _T_346 = _T_345 & io_exjump; // @[preBranch.scala 49:55]
  wire  _T_348 = _T_346 & _T_340; // @[preBranch.scala 49:67]
  wire  _T_350 = _T_348 & _T_52; // @[preBranch.scala 49:82]
  wire  _GEN_31 = _T_350 | vList_15; // @[Reg.scala 28:19]
  wire  _T_359 = io_ifpc == pcList_0; // @[preBranch.scala 58:29]
  wire  hitIfList_0 = _T_359 & vList_0; // @[preBranch.scala 58:43]
  wire  _T_361 = io_ifpc == pcList_1; // @[preBranch.scala 58:29]
  wire  hitIfList_1 = _T_361 & vList_1; // @[preBranch.scala 58:43]
  wire  _T_363 = io_ifpc == pcList_2; // @[preBranch.scala 58:29]
  wire  hitIfList_2 = _T_363 & vList_2; // @[preBranch.scala 58:43]
  wire  _T_365 = io_ifpc == pcList_3; // @[preBranch.scala 58:29]
  wire  hitIfList_3 = _T_365 & vList_3; // @[preBranch.scala 58:43]
  wire  _T_367 = io_ifpc == pcList_4; // @[preBranch.scala 58:29]
  wire  hitIfList_4 = _T_367 & vList_4; // @[preBranch.scala 58:43]
  wire  _T_369 = io_ifpc == pcList_5; // @[preBranch.scala 58:29]
  wire  hitIfList_5 = _T_369 & vList_5; // @[preBranch.scala 58:43]
  wire  _T_371 = io_ifpc == pcList_6; // @[preBranch.scala 58:29]
  wire  hitIfList_6 = _T_371 & vList_6; // @[preBranch.scala 58:43]
  wire  _T_373 = io_ifpc == pcList_7; // @[preBranch.scala 58:29]
  wire  hitIfList_7 = _T_373 & vList_7; // @[preBranch.scala 58:43]
  wire  _T_375 = io_ifpc == pcList_8; // @[preBranch.scala 58:29]
  wire  hitIfList_8 = _T_375 & vList_8; // @[preBranch.scala 58:43]
  wire  _T_377 = io_ifpc == pcList_9; // @[preBranch.scala 58:29]
  wire  hitIfList_9 = _T_377 & vList_9; // @[preBranch.scala 58:43]
  wire  _T_379 = io_ifpc == pcList_10; // @[preBranch.scala 58:29]
  wire  hitIfList_10 = _T_379 & vList_10; // @[preBranch.scala 58:43]
  wire  _T_381 = io_ifpc == pcList_11; // @[preBranch.scala 58:29]
  wire  hitIfList_11 = _T_381 & vList_11; // @[preBranch.scala 58:43]
  wire  _T_383 = io_ifpc == pcList_12; // @[preBranch.scala 58:29]
  wire  hitIfList_12 = _T_383 & vList_12; // @[preBranch.scala 58:43]
  wire  _T_385 = io_ifpc == pcList_13; // @[preBranch.scala 58:29]
  wire  hitIfList_13 = _T_385 & vList_13; // @[preBranch.scala 58:43]
  wire  _T_387 = io_ifpc == pcList_14; // @[preBranch.scala 58:29]
  wire  hitIfList_14 = _T_387 & vList_14; // @[preBranch.scala 58:43]
  wire  _T_389 = io_ifpc == pcList_15; // @[preBranch.scala 58:29]
  wire  hitIfList_15 = _T_389 & vList_15; // @[preBranch.scala 58:43]
  wire  _T_392 = hitIfList_0 | hitIfList_1; // @[preBranch.scala 61:55]
  wire  _T_393 = _T_392 | hitIfList_2; // @[preBranch.scala 61:55]
  wire  _T_394 = _T_393 | hitIfList_3; // @[preBranch.scala 61:55]
  wire  _T_395 = _T_394 | hitIfList_4; // @[preBranch.scala 61:55]
  wire  _T_396 = _T_395 | hitIfList_5; // @[preBranch.scala 61:55]
  wire  _T_397 = _T_396 | hitIfList_6; // @[preBranch.scala 61:55]
  wire  _T_398 = _T_397 | hitIfList_7; // @[preBranch.scala 61:55]
  wire  _T_399 = _T_398 | hitIfList_8; // @[preBranch.scala 61:55]
  wire  _T_400 = _T_399 | hitIfList_9; // @[preBranch.scala 61:55]
  wire  _T_401 = _T_400 | hitIfList_10; // @[preBranch.scala 61:55]
  wire  _T_402 = _T_401 | hitIfList_11; // @[preBranch.scala 61:55]
  wire  _T_403 = _T_402 | hitIfList_12; // @[preBranch.scala 61:55]
  wire  _T_404 = _T_403 | hitIfList_13; // @[preBranch.scala 61:55]
  wire  _T_405 = _T_404 | hitIfList_14; // @[preBranch.scala 61:55]
  wire  hitif = _T_405 | hitIfList_15; // @[preBranch.scala 61:55]
  wire  _T_406 = ~hitif; // @[preBranch.scala 67:5]
  wire  _T_407 = hitIfList_0 & precelList_0_io_valid; // @[Mux.scala 27:72]
  wire  _T_408 = hitIfList_1 & precelList_1_io_valid; // @[Mux.scala 27:72]
  wire  _T_409 = hitIfList_2 & precelList_2_io_valid; // @[Mux.scala 27:72]
  wire  _T_410 = hitIfList_3 & precelList_3_io_valid; // @[Mux.scala 27:72]
  wire  _T_411 = hitIfList_4 & precelList_4_io_valid; // @[Mux.scala 27:72]
  wire  _T_412 = hitIfList_5 & precelList_5_io_valid; // @[Mux.scala 27:72]
  wire  _T_413 = hitIfList_6 & precelList_6_io_valid; // @[Mux.scala 27:72]
  wire  _T_414 = hitIfList_7 & precelList_7_io_valid; // @[Mux.scala 27:72]
  wire  _T_415 = hitIfList_8 & precelList_8_io_valid; // @[Mux.scala 27:72]
  wire  _T_416 = hitIfList_9 & precelList_9_io_valid; // @[Mux.scala 27:72]
  wire  _T_417 = hitIfList_10 & precelList_10_io_valid; // @[Mux.scala 27:72]
  wire  _T_418 = hitIfList_11 & precelList_11_io_valid; // @[Mux.scala 27:72]
  wire  _T_419 = hitIfList_12 & precelList_12_io_valid; // @[Mux.scala 27:72]
  wire  _T_420 = hitIfList_13 & precelList_13_io_valid; // @[Mux.scala 27:72]
  wire  _T_421 = hitIfList_14 & precelList_14_io_valid; // @[Mux.scala 27:72]
  wire  _T_422 = hitIfList_15 & precelList_15_io_valid; // @[Mux.scala 27:72]
  wire  _T_423 = _T_407 | _T_408; // @[Mux.scala 27:72]
  wire  _T_424 = _T_423 | _T_409; // @[Mux.scala 27:72]
  wire  _T_425 = _T_424 | _T_410; // @[Mux.scala 27:72]
  wire  _T_426 = _T_425 | _T_411; // @[Mux.scala 27:72]
  wire  _T_427 = _T_426 | _T_412; // @[Mux.scala 27:72]
  wire  _T_428 = _T_427 | _T_413; // @[Mux.scala 27:72]
  wire  _T_429 = _T_428 | _T_414; // @[Mux.scala 27:72]
  wire  _T_430 = _T_429 | _T_415; // @[Mux.scala 27:72]
  wire  _T_431 = _T_430 | _T_416; // @[Mux.scala 27:72]
  wire  _T_432 = _T_431 | _T_417; // @[Mux.scala 27:72]
  wire  _T_433 = _T_432 | _T_418; // @[Mux.scala 27:72]
  wire  _T_434 = _T_433 | _T_419; // @[Mux.scala 27:72]
  wire  _T_435 = _T_434 | _T_420; // @[Mux.scala 27:72]
  wire  _T_436 = _T_435 | _T_421; // @[Mux.scala 27:72]
  wire  _T_437 = _T_436 | _T_422; // @[Mux.scala 27:72]
  wire [31:0] _T_441 = hitIfList_0 ? precelList_0_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_442 = hitIfList_1 ? precelList_1_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_443 = hitIfList_2 ? precelList_2_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_444 = hitIfList_3 ? precelList_3_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_445 = hitIfList_4 ? precelList_4_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_446 = hitIfList_5 ? precelList_5_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_447 = hitIfList_6 ? precelList_6_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_448 = hitIfList_7 ? precelList_7_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_449 = hitIfList_8 ? precelList_8_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_450 = hitIfList_9 ? precelList_9_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_451 = hitIfList_10 ? precelList_10_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_452 = hitIfList_11 ? precelList_11_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_453 = hitIfList_12 ? precelList_12_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_454 = hitIfList_13 ? precelList_13_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_455 = hitIfList_14 ? precelList_14_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_456 = hitIfList_15 ? precelList_15_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_457 = _T_441 | _T_442; // @[Mux.scala 27:72]
  wire [31:0] _T_458 = _T_457 | _T_443; // @[Mux.scala 27:72]
  wire [31:0] _T_459 = _T_458 | _T_444; // @[Mux.scala 27:72]
  wire [31:0] _T_460 = _T_459 | _T_445; // @[Mux.scala 27:72]
  wire [31:0] _T_461 = _T_460 | _T_446; // @[Mux.scala 27:72]
  wire [31:0] _T_462 = _T_461 | _T_447; // @[Mux.scala 27:72]
  wire [31:0] _T_463 = _T_462 | _T_448; // @[Mux.scala 27:72]
  wire [31:0] _T_464 = _T_463 | _T_449; // @[Mux.scala 27:72]
  wire [31:0] _T_465 = _T_464 | _T_450; // @[Mux.scala 27:72]
  wire [31:0] _T_466 = _T_465 | _T_451; // @[Mux.scala 27:72]
  wire [31:0] _T_467 = _T_466 | _T_452; // @[Mux.scala 27:72]
  wire [31:0] _T_468 = _T_467 | _T_453; // @[Mux.scala 27:72]
  wire [31:0] _T_469 = _T_468 | _T_454; // @[Mux.scala 27:72]
  wire [31:0] _T_470 = _T_469 | _T_455; // @[Mux.scala 27:72]
  wire [31:0] _T_471 = _T_470 | _T_456; // @[Mux.scala 27:72]
  preCell precelList_0 ( // @[preBranch.scala 30:45]
    .clock(precelList_0_clock),
    .reset(precelList_0_reset),
    .io_cen(precelList_0_io_cen),
    .io_jump(precelList_0_io_jump),
    .io_dnpcIn(precelList_0_io_dnpcIn),
    .io_dnpcOut(precelList_0_io_dnpcOut),
    .io_valid(precelList_0_io_valid)
  );
  preCell precelList_1 ( // @[preBranch.scala 30:45]
    .clock(precelList_1_clock),
    .reset(precelList_1_reset),
    .io_cen(precelList_1_io_cen),
    .io_jump(precelList_1_io_jump),
    .io_dnpcIn(precelList_1_io_dnpcIn),
    .io_dnpcOut(precelList_1_io_dnpcOut),
    .io_valid(precelList_1_io_valid)
  );
  preCell precelList_2 ( // @[preBranch.scala 30:45]
    .clock(precelList_2_clock),
    .reset(precelList_2_reset),
    .io_cen(precelList_2_io_cen),
    .io_jump(precelList_2_io_jump),
    .io_dnpcIn(precelList_2_io_dnpcIn),
    .io_dnpcOut(precelList_2_io_dnpcOut),
    .io_valid(precelList_2_io_valid)
  );
  preCell precelList_3 ( // @[preBranch.scala 30:45]
    .clock(precelList_3_clock),
    .reset(precelList_3_reset),
    .io_cen(precelList_3_io_cen),
    .io_jump(precelList_3_io_jump),
    .io_dnpcIn(precelList_3_io_dnpcIn),
    .io_dnpcOut(precelList_3_io_dnpcOut),
    .io_valid(precelList_3_io_valid)
  );
  preCell precelList_4 ( // @[preBranch.scala 30:45]
    .clock(precelList_4_clock),
    .reset(precelList_4_reset),
    .io_cen(precelList_4_io_cen),
    .io_jump(precelList_4_io_jump),
    .io_dnpcIn(precelList_4_io_dnpcIn),
    .io_dnpcOut(precelList_4_io_dnpcOut),
    .io_valid(precelList_4_io_valid)
  );
  preCell precelList_5 ( // @[preBranch.scala 30:45]
    .clock(precelList_5_clock),
    .reset(precelList_5_reset),
    .io_cen(precelList_5_io_cen),
    .io_jump(precelList_5_io_jump),
    .io_dnpcIn(precelList_5_io_dnpcIn),
    .io_dnpcOut(precelList_5_io_dnpcOut),
    .io_valid(precelList_5_io_valid)
  );
  preCell precelList_6 ( // @[preBranch.scala 30:45]
    .clock(precelList_6_clock),
    .reset(precelList_6_reset),
    .io_cen(precelList_6_io_cen),
    .io_jump(precelList_6_io_jump),
    .io_dnpcIn(precelList_6_io_dnpcIn),
    .io_dnpcOut(precelList_6_io_dnpcOut),
    .io_valid(precelList_6_io_valid)
  );
  preCell precelList_7 ( // @[preBranch.scala 30:45]
    .clock(precelList_7_clock),
    .reset(precelList_7_reset),
    .io_cen(precelList_7_io_cen),
    .io_jump(precelList_7_io_jump),
    .io_dnpcIn(precelList_7_io_dnpcIn),
    .io_dnpcOut(precelList_7_io_dnpcOut),
    .io_valid(precelList_7_io_valid)
  );
  preCell precelList_8 ( // @[preBranch.scala 30:45]
    .clock(precelList_8_clock),
    .reset(precelList_8_reset),
    .io_cen(precelList_8_io_cen),
    .io_jump(precelList_8_io_jump),
    .io_dnpcIn(precelList_8_io_dnpcIn),
    .io_dnpcOut(precelList_8_io_dnpcOut),
    .io_valid(precelList_8_io_valid)
  );
  preCell precelList_9 ( // @[preBranch.scala 30:45]
    .clock(precelList_9_clock),
    .reset(precelList_9_reset),
    .io_cen(precelList_9_io_cen),
    .io_jump(precelList_9_io_jump),
    .io_dnpcIn(precelList_9_io_dnpcIn),
    .io_dnpcOut(precelList_9_io_dnpcOut),
    .io_valid(precelList_9_io_valid)
  );
  preCell precelList_10 ( // @[preBranch.scala 30:45]
    .clock(precelList_10_clock),
    .reset(precelList_10_reset),
    .io_cen(precelList_10_io_cen),
    .io_jump(precelList_10_io_jump),
    .io_dnpcIn(precelList_10_io_dnpcIn),
    .io_dnpcOut(precelList_10_io_dnpcOut),
    .io_valid(precelList_10_io_valid)
  );
  preCell precelList_11 ( // @[preBranch.scala 30:45]
    .clock(precelList_11_clock),
    .reset(precelList_11_reset),
    .io_cen(precelList_11_io_cen),
    .io_jump(precelList_11_io_jump),
    .io_dnpcIn(precelList_11_io_dnpcIn),
    .io_dnpcOut(precelList_11_io_dnpcOut),
    .io_valid(precelList_11_io_valid)
  );
  preCell precelList_12 ( // @[preBranch.scala 30:45]
    .clock(precelList_12_clock),
    .reset(precelList_12_reset),
    .io_cen(precelList_12_io_cen),
    .io_jump(precelList_12_io_jump),
    .io_dnpcIn(precelList_12_io_dnpcIn),
    .io_dnpcOut(precelList_12_io_dnpcOut),
    .io_valid(precelList_12_io_valid)
  );
  preCell precelList_13 ( // @[preBranch.scala 30:45]
    .clock(precelList_13_clock),
    .reset(precelList_13_reset),
    .io_cen(precelList_13_io_cen),
    .io_jump(precelList_13_io_jump),
    .io_dnpcIn(precelList_13_io_dnpcIn),
    .io_dnpcOut(precelList_13_io_dnpcOut),
    .io_valid(precelList_13_io_valid)
  );
  preCell precelList_14 ( // @[preBranch.scala 30:45]
    .clock(precelList_14_clock),
    .reset(precelList_14_reset),
    .io_cen(precelList_14_io_cen),
    .io_jump(precelList_14_io_jump),
    .io_dnpcIn(precelList_14_io_dnpcIn),
    .io_dnpcOut(precelList_14_io_dnpcOut),
    .io_valid(precelList_14_io_valid)
  );
  preCell precelList_15 ( // @[preBranch.scala 30:45]
    .clock(precelList_15_clock),
    .reset(precelList_15_reset),
    .io_cen(precelList_15_io_cen),
    .io_jump(precelList_15_io_jump),
    .io_dnpcIn(precelList_15_io_dnpcIn),
    .io_dnpcOut(precelList_15_io_dnpcOut),
    .io_valid(precelList_15_io_valid)
  );
  assign io_ifdnpc = _T_406 ? 32'h0 : _T_471; // @[preBranch.scala 78:13]
  assign io_ifjump = _T_406 ? 1'h0 : _T_437; // @[preBranch.scala 66:13]
  assign precelList_0_clock = clock;
  assign precelList_0_reset = reset;
  assign precelList_0_io_cen = _T_57 & _T_52; // @[preBranch.scala 47:26]
  assign precelList_0_io_jump = io_exjump; // @[preBranch.scala 45:27]
  assign precelList_0_io_dnpcIn = io_exdpc; // @[preBranch.scala 46:29]
  assign precelList_1_clock = clock;
  assign precelList_1_reset = reset;
  assign precelList_1_io_cen = _T_76 & _T_52; // @[preBranch.scala 47:26]
  assign precelList_1_io_jump = io_exjump; // @[preBranch.scala 45:27]
  assign precelList_1_io_dnpcIn = io_exdpc; // @[preBranch.scala 46:29]
  assign precelList_2_clock = clock;
  assign precelList_2_reset = reset;
  assign precelList_2_io_cen = _T_95 & _T_52; // @[preBranch.scala 47:26]
  assign precelList_2_io_jump = io_exjump; // @[preBranch.scala 45:27]
  assign precelList_2_io_dnpcIn = io_exdpc; // @[preBranch.scala 46:29]
  assign precelList_3_clock = clock;
  assign precelList_3_reset = reset;
  assign precelList_3_io_cen = _T_114 & _T_52; // @[preBranch.scala 47:26]
  assign precelList_3_io_jump = io_exjump; // @[preBranch.scala 45:27]
  assign precelList_3_io_dnpcIn = io_exdpc; // @[preBranch.scala 46:29]
  assign precelList_4_clock = clock;
  assign precelList_4_reset = reset;
  assign precelList_4_io_cen = _T_133 & _T_52; // @[preBranch.scala 47:26]
  assign precelList_4_io_jump = io_exjump; // @[preBranch.scala 45:27]
  assign precelList_4_io_dnpcIn = io_exdpc; // @[preBranch.scala 46:29]
  assign precelList_5_clock = clock;
  assign precelList_5_reset = reset;
  assign precelList_5_io_cen = _T_152 & _T_52; // @[preBranch.scala 47:26]
  assign precelList_5_io_jump = io_exjump; // @[preBranch.scala 45:27]
  assign precelList_5_io_dnpcIn = io_exdpc; // @[preBranch.scala 46:29]
  assign precelList_6_clock = clock;
  assign precelList_6_reset = reset;
  assign precelList_6_io_cen = _T_171 & _T_52; // @[preBranch.scala 47:26]
  assign precelList_6_io_jump = io_exjump; // @[preBranch.scala 45:27]
  assign precelList_6_io_dnpcIn = io_exdpc; // @[preBranch.scala 46:29]
  assign precelList_7_clock = clock;
  assign precelList_7_reset = reset;
  assign precelList_7_io_cen = _T_190 & _T_52; // @[preBranch.scala 47:26]
  assign precelList_7_io_jump = io_exjump; // @[preBranch.scala 45:27]
  assign precelList_7_io_dnpcIn = io_exdpc; // @[preBranch.scala 46:29]
  assign precelList_8_clock = clock;
  assign precelList_8_reset = reset;
  assign precelList_8_io_cen = _T_209 & _T_52; // @[preBranch.scala 47:26]
  assign precelList_8_io_jump = io_exjump; // @[preBranch.scala 45:27]
  assign precelList_8_io_dnpcIn = io_exdpc; // @[preBranch.scala 46:29]
  assign precelList_9_clock = clock;
  assign precelList_9_reset = reset;
  assign precelList_9_io_cen = _T_228 & _T_52; // @[preBranch.scala 47:26]
  assign precelList_9_io_jump = io_exjump; // @[preBranch.scala 45:27]
  assign precelList_9_io_dnpcIn = io_exdpc; // @[preBranch.scala 46:29]
  assign precelList_10_clock = clock;
  assign precelList_10_reset = reset;
  assign precelList_10_io_cen = _T_247 & _T_52; // @[preBranch.scala 47:26]
  assign precelList_10_io_jump = io_exjump; // @[preBranch.scala 45:27]
  assign precelList_10_io_dnpcIn = io_exdpc; // @[preBranch.scala 46:29]
  assign precelList_11_clock = clock;
  assign precelList_11_reset = reset;
  assign precelList_11_io_cen = _T_266 & _T_52; // @[preBranch.scala 47:26]
  assign precelList_11_io_jump = io_exjump; // @[preBranch.scala 45:27]
  assign precelList_11_io_dnpcIn = io_exdpc; // @[preBranch.scala 46:29]
  assign precelList_12_clock = clock;
  assign precelList_12_reset = reset;
  assign precelList_12_io_cen = _T_285 & _T_52; // @[preBranch.scala 47:26]
  assign precelList_12_io_jump = io_exjump; // @[preBranch.scala 45:27]
  assign precelList_12_io_dnpcIn = io_exdpc; // @[preBranch.scala 46:29]
  assign precelList_13_clock = clock;
  assign precelList_13_reset = reset;
  assign precelList_13_io_cen = _T_304 & _T_52; // @[preBranch.scala 47:26]
  assign precelList_13_io_jump = io_exjump; // @[preBranch.scala 45:27]
  assign precelList_13_io_dnpcIn = io_exdpc; // @[preBranch.scala 46:29]
  assign precelList_14_clock = clock;
  assign precelList_14_reset = reset;
  assign precelList_14_io_cen = _T_323 & _T_52; // @[preBranch.scala 47:26]
  assign precelList_14_io_jump = io_exjump; // @[preBranch.scala 45:27]
  assign precelList_14_io_dnpcIn = io_exdpc; // @[preBranch.scala 46:29]
  assign precelList_15_clock = clock;
  assign precelList_15_reset = reset;
  assign precelList_15_io_cen = _T_342 & _T_52; // @[preBranch.scala 47:26]
  assign precelList_15_io_jump = io_exjump; // @[preBranch.scala 45:27]
  assign precelList_15_io_dnpcIn = io_exdpc; // @[preBranch.scala 46:29]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pcList_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  vList_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  pcList_1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  vList_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  pcList_2 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  vList_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  pcList_3 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  vList_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  pcList_4 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  vList_4 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  pcList_5 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  vList_5 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  pcList_6 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  vList_6 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  pcList_7 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  vList_7 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  pcList_8 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  vList_8 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  pcList_9 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  vList_9 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  pcList_10 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  vList_10 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  pcList_11 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  vList_11 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  pcList_12 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  vList_12 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  pcList_13 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  vList_13 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  pcList_14 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  vList_14 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  pcList_15 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  vList_15 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  cnt = _RAND_32[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pcList_0 <= 32'h0;
    end else if (_T_65) begin
      pcList_0 <= io_expc;
    end
    if (reset) begin
      vList_0 <= 1'h0;
    end else begin
      vList_0 <= _GEN_1;
    end
    if (reset) begin
      pcList_1 <= 32'h0;
    end else if (_T_84) begin
      pcList_1 <= io_expc;
    end
    if (reset) begin
      vList_1 <= 1'h0;
    end else begin
      vList_1 <= _GEN_3;
    end
    if (reset) begin
      pcList_2 <= 32'h0;
    end else if (_T_103) begin
      pcList_2 <= io_expc;
    end
    if (reset) begin
      vList_2 <= 1'h0;
    end else begin
      vList_2 <= _GEN_5;
    end
    if (reset) begin
      pcList_3 <= 32'h0;
    end else if (_T_122) begin
      pcList_3 <= io_expc;
    end
    if (reset) begin
      vList_3 <= 1'h0;
    end else begin
      vList_3 <= _GEN_7;
    end
    if (reset) begin
      pcList_4 <= 32'h0;
    end else if (_T_141) begin
      pcList_4 <= io_expc;
    end
    if (reset) begin
      vList_4 <= 1'h0;
    end else begin
      vList_4 <= _GEN_9;
    end
    if (reset) begin
      pcList_5 <= 32'h0;
    end else if (_T_160) begin
      pcList_5 <= io_expc;
    end
    if (reset) begin
      vList_5 <= 1'h0;
    end else begin
      vList_5 <= _GEN_11;
    end
    if (reset) begin
      pcList_6 <= 32'h0;
    end else if (_T_179) begin
      pcList_6 <= io_expc;
    end
    if (reset) begin
      vList_6 <= 1'h0;
    end else begin
      vList_6 <= _GEN_13;
    end
    if (reset) begin
      pcList_7 <= 32'h0;
    end else if (_T_198) begin
      pcList_7 <= io_expc;
    end
    if (reset) begin
      vList_7 <= 1'h0;
    end else begin
      vList_7 <= _GEN_15;
    end
    if (reset) begin
      pcList_8 <= 32'h0;
    end else if (_T_217) begin
      pcList_8 <= io_expc;
    end
    if (reset) begin
      vList_8 <= 1'h0;
    end else begin
      vList_8 <= _GEN_17;
    end
    if (reset) begin
      pcList_9 <= 32'h0;
    end else if (_T_236) begin
      pcList_9 <= io_expc;
    end
    if (reset) begin
      vList_9 <= 1'h0;
    end else begin
      vList_9 <= _GEN_19;
    end
    if (reset) begin
      pcList_10 <= 32'h0;
    end else if (_T_255) begin
      pcList_10 <= io_expc;
    end
    if (reset) begin
      vList_10 <= 1'h0;
    end else begin
      vList_10 <= _GEN_21;
    end
    if (reset) begin
      pcList_11 <= 32'h0;
    end else if (_T_274) begin
      pcList_11 <= io_expc;
    end
    if (reset) begin
      vList_11 <= 1'h0;
    end else begin
      vList_11 <= _GEN_23;
    end
    if (reset) begin
      pcList_12 <= 32'h0;
    end else if (_T_293) begin
      pcList_12 <= io_expc;
    end
    if (reset) begin
      vList_12 <= 1'h0;
    end else begin
      vList_12 <= _GEN_25;
    end
    if (reset) begin
      pcList_13 <= 32'h0;
    end else if (_T_312) begin
      pcList_13 <= io_expc;
    end
    if (reset) begin
      vList_13 <= 1'h0;
    end else begin
      vList_13 <= _GEN_27;
    end
    if (reset) begin
      pcList_14 <= 32'h0;
    end else if (_T_331) begin
      pcList_14 <= io_expc;
    end
    if (reset) begin
      vList_14 <= 1'h0;
    end else begin
      vList_14 <= _GEN_29;
    end
    if (reset) begin
      pcList_15 <= 32'h0;
    end else if (_T_350) begin
      pcList_15 <= io_expc;
    end
    if (reset) begin
      vList_15 <= 1'h0;
    end else begin
      vList_15 <= _GEN_31;
    end
    if (reset) begin
      cnt <= 4'h0;
    end else if (_T_53) begin
      cnt <= _T_49;
    end
  end
endmodule
module memVGen(
  input  [31:0] io_inst,
  output        io_valid
);
  wire [31:0] _T = io_inst & 32'h707f; // @[memVGen.scala 21:45]
  wire  _T_1 = 32'h3023 == _T; // @[memVGen.scala 21:45]
  wire  _T_3 = 32'h2023 == _T; // @[memVGen.scala 21:45]
  wire  _T_5 = 32'h23 == _T; // @[memVGen.scala 21:45]
  wire  _T_7 = 32'h1023 == _T; // @[memVGen.scala 21:45]
  wire  _T_9 = 32'h3003 == _T; // @[memVGen.scala 27:27]
  wire  _T_11 = 32'h4003 == _T; // @[memVGen.scala 28:27]
  wire  _T_13 = 32'h1003 == _T; // @[memVGen.scala 29:27]
  wire  _T_15 = 32'h2003 == _T; // @[memVGen.scala 30:27]
  wire  _T_19 = 32'h5003 == _T; // @[memVGen.scala 32:27]
  wire  _T_21 = 32'h3 == _T; // @[memVGen.scala 33:27]
  wire  _T_23 = 32'h6003 == _T; // @[memVGen.scala 34:27]
  wire  _T_25 = _T_21 | _T_23; // @[Mux.scala 98:16]
  wire  _T_26 = _T_19 | _T_25; // @[Mux.scala 98:16]
  wire  _T_27 = _T_9 | _T_26; // @[Mux.scala 98:16]
  wire  _T_28 = _T_15 | _T_27; // @[Mux.scala 98:16]
  wire  _T_29 = _T_13 | _T_28; // @[Mux.scala 98:16]
  wire  _T_30 = _T_11 | _T_29; // @[Mux.scala 98:16]
  wire  _T_31 = _T_9 | _T_30; // @[Mux.scala 98:16]
  wire  _T_32 = _T_7 | _T_31; // @[Mux.scala 98:16]
  wire  _T_33 = _T_5 | _T_32; // @[Mux.scala 98:16]
  wire  _T_34 = _T_3 | _T_33; // @[Mux.scala 98:16]
  assign io_valid = _T_1 | _T_34; // @[memVGen.scala 37:12]
endmodule
module ALUCtrl(
  input  [31:0] io_inst,
  output [4:0]  io_ALUCtrl
);
  wire [31:0] _T = io_inst & 32'h707f; // @[ALUCtrl.scala 75:49]
  wire  _T_1 = 32'h3023 == _T; // @[ALUCtrl.scala 75:49]
  wire  _T_3 = 32'h2023 == _T; // @[ALUCtrl.scala 75:49]
  wire  _T_5 = 32'h23 == _T; // @[ALUCtrl.scala 75:49]
  wire  _T_7 = 32'h1023 == _T; // @[ALUCtrl.scala 75:49]
  wire [31:0] _T_8 = io_inst & 32'h7f; // @[ALUCtrl.scala 80:31]
  wire  _T_9 = 32'h17 == _T_8; // @[ALUCtrl.scala 80:31]
  wire  _T_11 = 32'h37 == _T_8; // @[ALUCtrl.scala 81:31]
  wire  _T_13 = 32'h13 == _T; // @[ALUCtrl.scala 82:31]
  wire  _T_15 = 32'h67 == _T; // @[ALUCtrl.scala 83:31]
  wire  _T_17 = 32'h3003 == _T; // @[ALUCtrl.scala 84:31]
  wire  _T_19 = 32'h4003 == _T; // @[ALUCtrl.scala 85:31]
  wire  _T_21 = 32'h3013 == _T; // @[ALUCtrl.scala 86:31]
  wire [31:0] _T_22 = io_inst & 32'hfe00707f; // @[ALUCtrl.scala 87:31]
  wire  _T_23 = 32'h501b == _T_22; // @[ALUCtrl.scala 87:31]
  wire [31:0] _T_24 = io_inst & 32'hfc00707f; // @[ALUCtrl.scala 88:31]
  wire  _T_25 = 32'h1013 == _T_24; // @[ALUCtrl.scala 88:31]
  wire  _T_27 = 32'h7013 == _T; // @[ALUCtrl.scala 89:31]
  wire  _T_29 = 32'h4013 == _T; // @[ALUCtrl.scala 90:31]
  wire  _T_31 = 32'h1b == _T; // @[ALUCtrl.scala 91:31]
  wire  _T_33 = 32'h5013 == _T_24; // @[ALUCtrl.scala 92:31]
  wire  _T_35 = 32'h101b == _T_22; // @[ALUCtrl.scala 93:31]
  wire  _T_37 = 32'h4000501b == _T_22; // @[ALUCtrl.scala 94:31]
  wire  _T_39 = 32'h40005013 == _T_24; // @[ALUCtrl.scala 95:31]
  wire  _T_41 = 32'h1003 == _T; // @[ALUCtrl.scala 96:31]
  wire  _T_43 = 32'h2003 == _T; // @[ALUCtrl.scala 97:31]
  wire  _T_47 = 32'h5003 == _T; // @[ALUCtrl.scala 99:31]
  wire  _T_49 = 32'h6003 == _T; // @[ALUCtrl.scala 100:31]
  wire  _T_51 = 32'h3 == _T; // @[ALUCtrl.scala 101:31]
  wire  _T_53 = 32'h6013 == _T; // @[ALUCtrl.scala 102:31]
  wire  _T_55 = 32'h3033 == _T_22; // @[ALUCtrl.scala 103:31]
  wire  _T_57 = 32'h3b == _T_22; // @[ALUCtrl.scala 104:31]
  wire  _T_59 = 32'h4000003b == _T_22; // @[ALUCtrl.scala 105:31]
  wire  _T_61 = 32'h7033 == _T_22; // @[ALUCtrl.scala 106:31]
  wire  _T_63 = 32'h33 == _T_22; // @[ALUCtrl.scala 107:31]
  wire  _T_65 = 32'h200503b == _T_22; // @[ALUCtrl.scala 108:31]
  wire  _T_67 = 32'h200703b == _T_22; // @[ALUCtrl.scala 109:31]
  wire  _T_69 = 32'h40000033 == _T_22; // @[ALUCtrl.scala 110:31]
  wire  _T_71 = 32'h200003b == _T_22; // @[ALUCtrl.scala 111:31]
  wire  _T_73 = 32'h200603b == _T_22; // @[ALUCtrl.scala 112:31]
  wire  _T_75 = 32'h200403b == _T_22; // @[ALUCtrl.scala 113:31]
  wire  _T_77 = 32'h2000033 == _T_22; // @[ALUCtrl.scala 114:31]
  wire  _T_79 = 32'h6033 == _T_22; // @[ALUCtrl.scala 115:31]
  wire  _T_81 = 32'h103b == _T_22; // @[ALUCtrl.scala 116:31]
  wire  _T_83 = 32'h4000503b == _T_22; // @[ALUCtrl.scala 117:31]
  wire  _T_85 = 32'h503b == _T_22; // @[ALUCtrl.scala 118:31]
  wire  _T_87 = 32'h2033 == _T_22; // @[ALUCtrl.scala 119:31]
  wire  _T_89 = 32'h2005033 == _T_22; // @[ALUCtrl.scala 120:31]
  wire  _T_91 = 32'h4033 == _T_22; // @[ALUCtrl.scala 121:31]
  wire  _T_93 = 32'h2006033 == _T_22; // @[ALUCtrl.scala 122:31]
  wire  _T_95 = 32'h2004033 == _T_22; // @[ALUCtrl.scala 123:31]
  wire  _T_97 = 32'h1033 == _T_22; // @[ALUCtrl.scala 124:31]
  wire  _T_99 = 32'h63 == _T; // @[ALUCtrl.scala 125:31]
  wire  _T_101 = 32'h6063 == _T; // @[ALUCtrl.scala 126:31]
  wire  _T_103 = 32'h7063 == _T; // @[ALUCtrl.scala 127:31]
  wire  _T_105 = 32'h4063 == _T; // @[ALUCtrl.scala 128:31]
  wire  _T_107 = 32'h5063 == _T; // @[ALUCtrl.scala 129:31]
  wire  _T_109 = 32'h1063 == _T; // @[ALUCtrl.scala 130:31]
  wire  _T_111 = 32'h2007033 == _T_22; // @[ALUCtrl.scala 131:31]
  wire  _T_113 = 32'h5033 == _T_22; // @[ALUCtrl.scala 132:31]
  wire [4:0] _T_114 = _T_113 ? 5'h8 : 5'h1f; // @[Mux.scala 98:16]
  wire [4:0] _T_115 = _T_111 ? 5'h1d : _T_114; // @[Mux.scala 98:16]
  wire [4:0] _T_116 = _T_109 ? 5'hb : _T_115; // @[Mux.scala 98:16]
  wire [4:0] _T_117 = _T_107 ? 5'h1c : _T_116; // @[Mux.scala 98:16]
  wire [4:0] _T_118 = _T_105 ? 5'h5 : _T_117; // @[Mux.scala 98:16]
  wire [4:0] _T_119 = _T_103 ? 5'h1b : _T_118; // @[Mux.scala 98:16]
  wire [4:0] _T_120 = _T_101 ? 5'h7 : _T_119; // @[Mux.scala 98:16]
  wire [4:0] _T_121 = _T_99 ? 5'h1a : _T_120; // @[Mux.scala 98:16]
  wire [4:0] _T_122 = _T_97 ? 5'h6 : _T_121; // @[Mux.scala 98:16]
  wire [4:0] _T_123 = _T_95 ? 5'h19 : _T_122; // @[Mux.scala 98:16]
  wire [4:0] _T_124 = _T_93 ? 5'h18 : _T_123; // @[Mux.scala 98:16]
  wire [4:0] _T_125 = _T_91 ? 5'h4 : _T_124; // @[Mux.scala 98:16]
  wire [4:0] _T_126 = _T_89 ? 5'h17 : _T_125; // @[Mux.scala 98:16]
  wire [4:0] _T_127 = _T_87 ? 5'h5 : _T_126; // @[Mux.scala 98:16]
  wire [4:0] _T_128 = _T_85 ? 5'hc : _T_127; // @[Mux.scala 98:16]
  wire [4:0] _T_129 = _T_83 ? 5'hf : _T_128; // @[Mux.scala 98:16]
  wire [4:0] _T_130 = _T_81 ? 5'he : _T_129; // @[Mux.scala 98:16]
  wire [4:0] _T_131 = _T_79 ? 5'h3 : _T_130; // @[Mux.scala 98:16]
  wire [4:0] _T_132 = _T_77 ? 5'h16 : _T_131; // @[Mux.scala 98:16]
  wire [4:0] _T_133 = _T_75 ? 5'h15 : _T_132; // @[Mux.scala 98:16]
  wire [4:0] _T_134 = _T_73 ? 5'h14 : _T_133; // @[Mux.scala 98:16]
  wire [4:0] _T_135 = _T_71 ? 5'h13 : _T_134; // @[Mux.scala 98:16]
  wire [4:0] _T_136 = _T_69 ? 5'h1 : _T_135; // @[Mux.scala 98:16]
  wire [4:0] _T_137 = _T_67 ? 5'h12 : _T_136; // @[Mux.scala 98:16]
  wire [4:0] _T_138 = _T_65 ? 5'h11 : _T_137; // @[Mux.scala 98:16]
  wire [4:0] _T_139 = _T_63 ? 5'h0 : _T_138; // @[Mux.scala 98:16]
  wire [4:0] _T_140 = _T_61 ? 5'h2 : _T_139; // @[Mux.scala 98:16]
  wire [4:0] _T_141 = _T_59 ? 5'h10 : _T_140; // @[Mux.scala 98:16]
  wire [4:0] _T_142 = _T_57 ? 5'hd : _T_141; // @[Mux.scala 98:16]
  wire [4:0] _T_143 = _T_55 ? 5'h7 : _T_142; // @[Mux.scala 98:16]
  wire [4:0] _T_144 = _T_53 ? 5'h3 : _T_143; // @[Mux.scala 98:16]
  wire [4:0] _T_145 = _T_51 ? 5'h0 : _T_144; // @[Mux.scala 98:16]
  wire [4:0] _T_146 = _T_49 ? 5'h0 : _T_145; // @[Mux.scala 98:16]
  wire [4:0] _T_147 = _T_47 ? 5'h0 : _T_146; // @[Mux.scala 98:16]
  wire [4:0] _T_148 = _T_17 ? 5'h0 : _T_147; // @[Mux.scala 98:16]
  wire [4:0] _T_149 = _T_43 ? 5'h0 : _T_148; // @[Mux.scala 98:16]
  wire [4:0] _T_150 = _T_41 ? 5'h0 : _T_149; // @[Mux.scala 98:16]
  wire [4:0] _T_151 = _T_39 ? 5'h9 : _T_150; // @[Mux.scala 98:16]
  wire [4:0] _T_152 = _T_37 ? 5'hf : _T_151; // @[Mux.scala 98:16]
  wire [4:0] _T_153 = _T_35 ? 5'he : _T_152; // @[Mux.scala 98:16]
  wire [4:0] _T_154 = _T_33 ? 5'h8 : _T_153; // @[Mux.scala 98:16]
  wire [4:0] _T_155 = _T_31 ? 5'hd : _T_154; // @[Mux.scala 98:16]
  wire [4:0] _T_156 = _T_29 ? 5'h4 : _T_155; // @[Mux.scala 98:16]
  wire [4:0] _T_157 = _T_27 ? 5'h2 : _T_156; // @[Mux.scala 98:16]
  wire [4:0] _T_158 = _T_25 ? 5'h6 : _T_157; // @[Mux.scala 98:16]
  wire [4:0] _T_159 = _T_23 ? 5'hc : _T_158; // @[Mux.scala 98:16]
  wire [4:0] _T_160 = _T_21 ? 5'h7 : _T_159; // @[Mux.scala 98:16]
  wire [4:0] _T_161 = _T_19 ? 5'h0 : _T_160; // @[Mux.scala 98:16]
  wire [4:0] _T_162 = _T_17 ? 5'h0 : _T_161; // @[Mux.scala 98:16]
  wire [4:0] _T_163 = _T_15 ? 5'h1f : _T_162; // @[Mux.scala 98:16]
  wire [4:0] _T_164 = _T_13 ? 5'h0 : _T_163; // @[Mux.scala 98:16]
  wire [4:0] _T_165 = _T_11 ? 5'ha : _T_164; // @[Mux.scala 98:16]
  wire [4:0] _T_166 = _T_9 ? 5'h0 : _T_165; // @[Mux.scala 98:16]
  wire [4:0] _T_167 = _T_7 ? 5'h0 : _T_166; // @[Mux.scala 98:16]
  wire [4:0] _T_168 = _T_5 ? 5'h0 : _T_167; // @[Mux.scala 98:16]
  wire [4:0] _T_169 = _T_3 ? 5'h0 : _T_168; // @[Mux.scala 98:16]
  assign io_ALUCtrl = _T_1 ? 5'h0 : _T_169; // @[ALUCtrl.scala 135:14]
endmodule
module ALUSrcGen(
  input  [31:0] io_inst,
  output [1:0]  io_AluSrc1,
  output [1:0]  io_AluSrc2
);
  wire [31:0] _T = io_inst & 32'hfe00707f; // @[ALUSrcGen.scala 67:49]
  wire  _T_1 = 32'h4033 == _T; // @[ALUSrcGen.scala 67:49]
  wire [31:0] _T_2 = io_inst & 32'h707f; // @[ALUSrcGen.scala 65:49]
  wire  _T_3 = 32'h3023 == _T_2; // @[ALUSrcGen.scala 65:49]
  wire [31:0] _T_4 = io_inst & 32'hfc00707f; // @[ALUSrcGen.scala 64:49]
  wire  _T_5 = 32'h1013 == _T_4; // @[ALUSrcGen.scala 64:49]
  wire  _T_7 = 32'h503b == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_9 = 32'h6063 == _T_2; // @[ALUSrcGen.scala 66:49]
  wire  _T_11 = 32'h1003 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire  _T_13 = 32'h2004033 == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_15 = 32'h4013 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire  _T_17 = 32'h2006033 == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_19 = 32'h200403b == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_21 = 32'h3033 == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_23 = 32'h6013 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire  _T_25 = 32'h5033 == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_27 = 32'h5063 == _T_2; // @[ALUSrcGen.scala 66:49]
  wire  _T_29 = 32'h6033 == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_31 = 32'h4000503b == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_33 = 32'h7013 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire  _T_35 = 32'h33 == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_37 = 32'h103b == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_39 = 32'h2000033 == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_41 = 32'h2005033 == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_43 = 32'h2033 == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_45 = 32'h4003 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire  _T_47 = 32'h3 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire  _T_49 = 32'h2023 == _T_2; // @[ALUSrcGen.scala 65:49]
  wire  _T_51 = 32'h200703b == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_53 = 32'h1063 == _T_2; // @[ALUSrcGen.scala 66:49]
  wire  _T_55 = 32'h1b == _T_2; // @[ALUSrcGen.scala 64:49]
  wire  _T_57 = 32'h4063 == _T_2; // @[ALUSrcGen.scala 66:49]
  wire  _T_59 = 32'h40005013 == _T_4; // @[ALUSrcGen.scala 64:49]
  wire  _T_61 = 32'h200603b == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_63 = 32'h63 == _T_2; // @[ALUSrcGen.scala 66:49]
  wire  _T_65 = 32'h3003 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire  _T_67 = 32'h3b == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_69 = 32'h4000501b == _T; // @[ALUSrcGen.scala 64:49]
  wire  _T_71 = 32'h7033 == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_73 = 32'h200003b == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_75 = 32'h67 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire  _T_77 = 32'h2007033 == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_79 = 32'h5013 == _T_4; // @[ALUSrcGen.scala 64:49]
  wire  _T_81 = 32'h4000003b == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_83 = 32'h200503b == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_85 = 32'h23 == _T_2; // @[ALUSrcGen.scala 65:49]
  wire  _T_87 = 32'h40000033 == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_89 = 32'h501b == _T; // @[ALUSrcGen.scala 64:49]
  wire  _T_91 = 32'h5003 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire  _T_93 = 32'h6003 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire  _T_95 = 32'h2003 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire  _T_97 = 32'h101b == _T; // @[ALUSrcGen.scala 64:49]
  wire  _T_99 = 32'h1023 == _T_2; // @[ALUSrcGen.scala 65:49]
  wire  _T_101 = 32'h13 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire  _T_103 = 32'h7063 == _T_2; // @[ALUSrcGen.scala 66:49]
  wire  _T_105 = 32'h1033 == _T; // @[ALUSrcGen.scala 67:49]
  wire  _T_107 = 32'h3013 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire [31:0] _T_108 = io_inst & 32'h7f; // @[ALUSrcGen.scala 72:31]
  wire  _T_109 = 32'h17 == _T_108; // @[ALUSrcGen.scala 72:31]
  wire  _T_111 = 32'h37 == _T_108; // @[ALUSrcGen.scala 73:31]
  wire  _T_225 = _T_109 | _T_111; // @[Mux.scala 98:16]
  wire  _T_226 = _T_107 ? 1'h0 : _T_225; // @[Mux.scala 98:16]
  wire  _T_227 = _T_105 ? 1'h0 : _T_226; // @[Mux.scala 98:16]
  wire  _T_228 = _T_103 ? 1'h0 : _T_227; // @[Mux.scala 98:16]
  wire  _T_229 = _T_101 ? 1'h0 : _T_228; // @[Mux.scala 98:16]
  wire  _T_230 = _T_99 ? 1'h0 : _T_229; // @[Mux.scala 98:16]
  wire  _T_231 = _T_97 ? 1'h0 : _T_230; // @[Mux.scala 98:16]
  wire  _T_232 = _T_95 ? 1'h0 : _T_231; // @[Mux.scala 98:16]
  wire  _T_233 = _T_93 ? 1'h0 : _T_232; // @[Mux.scala 98:16]
  wire  _T_234 = _T_91 ? 1'h0 : _T_233; // @[Mux.scala 98:16]
  wire  _T_235 = _T_89 ? 1'h0 : _T_234; // @[Mux.scala 98:16]
  wire  _T_236 = _T_87 ? 1'h0 : _T_235; // @[Mux.scala 98:16]
  wire  _T_237 = _T_85 ? 1'h0 : _T_236; // @[Mux.scala 98:16]
  wire  _T_238 = _T_83 ? 1'h0 : _T_237; // @[Mux.scala 98:16]
  wire  _T_239 = _T_81 ? 1'h0 : _T_238; // @[Mux.scala 98:16]
  wire  _T_240 = _T_79 ? 1'h0 : _T_239; // @[Mux.scala 98:16]
  wire  _T_241 = _T_77 ? 1'h0 : _T_240; // @[Mux.scala 98:16]
  wire  _T_242 = _T_75 ? 1'h0 : _T_241; // @[Mux.scala 98:16]
  wire  _T_243 = _T_73 ? 1'h0 : _T_242; // @[Mux.scala 98:16]
  wire  _T_244 = _T_71 ? 1'h0 : _T_243; // @[Mux.scala 98:16]
  wire  _T_245 = _T_69 ? 1'h0 : _T_244; // @[Mux.scala 98:16]
  wire  _T_246 = _T_67 ? 1'h0 : _T_245; // @[Mux.scala 98:16]
  wire  _T_247 = _T_65 ? 1'h0 : _T_246; // @[Mux.scala 98:16]
  wire  _T_248 = _T_63 ? 1'h0 : _T_247; // @[Mux.scala 98:16]
  wire  _T_249 = _T_61 ? 1'h0 : _T_248; // @[Mux.scala 98:16]
  wire  _T_250 = _T_59 ? 1'h0 : _T_249; // @[Mux.scala 98:16]
  wire  _T_251 = _T_57 ? 1'h0 : _T_250; // @[Mux.scala 98:16]
  wire  _T_252 = _T_55 ? 1'h0 : _T_251; // @[Mux.scala 98:16]
  wire  _T_253 = _T_53 ? 1'h0 : _T_252; // @[Mux.scala 98:16]
  wire  _T_254 = _T_51 ? 1'h0 : _T_253; // @[Mux.scala 98:16]
  wire  _T_255 = _T_49 ? 1'h0 : _T_254; // @[Mux.scala 98:16]
  wire  _T_256 = _T_47 ? 1'h0 : _T_255; // @[Mux.scala 98:16]
  wire  _T_257 = _T_45 ? 1'h0 : _T_256; // @[Mux.scala 98:16]
  wire  _T_258 = _T_43 ? 1'h0 : _T_257; // @[Mux.scala 98:16]
  wire  _T_259 = _T_41 ? 1'h0 : _T_258; // @[Mux.scala 98:16]
  wire  _T_260 = _T_39 ? 1'h0 : _T_259; // @[Mux.scala 98:16]
  wire  _T_261 = _T_37 ? 1'h0 : _T_260; // @[Mux.scala 98:16]
  wire  _T_262 = _T_35 ? 1'h0 : _T_261; // @[Mux.scala 98:16]
  wire  _T_263 = _T_33 ? 1'h0 : _T_262; // @[Mux.scala 98:16]
  wire  _T_264 = _T_31 ? 1'h0 : _T_263; // @[Mux.scala 98:16]
  wire  _T_265 = _T_29 ? 1'h0 : _T_264; // @[Mux.scala 98:16]
  wire  _T_266 = _T_27 ? 1'h0 : _T_265; // @[Mux.scala 98:16]
  wire  _T_267 = _T_25 ? 1'h0 : _T_266; // @[Mux.scala 98:16]
  wire  _T_268 = _T_23 ? 1'h0 : _T_267; // @[Mux.scala 98:16]
  wire  _T_269 = _T_21 ? 1'h0 : _T_268; // @[Mux.scala 98:16]
  wire  _T_270 = _T_19 ? 1'h0 : _T_269; // @[Mux.scala 98:16]
  wire  _T_271 = _T_17 ? 1'h0 : _T_270; // @[Mux.scala 98:16]
  wire  _T_272 = _T_15 ? 1'h0 : _T_271; // @[Mux.scala 98:16]
  wire  _T_273 = _T_13 ? 1'h0 : _T_272; // @[Mux.scala 98:16]
  wire  _T_274 = _T_11 ? 1'h0 : _T_273; // @[Mux.scala 98:16]
  wire  _T_275 = _T_9 ? 1'h0 : _T_274; // @[Mux.scala 98:16]
  wire  _T_276 = _T_7 ? 1'h0 : _T_275; // @[Mux.scala 98:16]
  wire  _T_277 = _T_5 ? 1'h0 : _T_276; // @[Mux.scala 98:16]
  wire  _T_278 = _T_3 ? 1'h0 : _T_277; // @[Mux.scala 98:16]
  wire  _T_279 = _T_1 ? 1'h0 : _T_278; // @[Mux.scala 98:16]
  wire [1:0] _T_280 = _T_111 ? 2'h3 : 2'h0; // @[Mux.scala 98:16]
  wire [1:0] _T_281 = _T_109 ? 2'h2 : _T_280; // @[Mux.scala 98:16]
  wire [1:0] _T_282 = _T_107 ? 2'h1 : _T_281; // @[Mux.scala 98:16]
  wire [1:0] _T_283 = _T_105 ? 2'h0 : _T_282; // @[Mux.scala 98:16]
  wire [1:0] _T_284 = _T_103 ? 2'h0 : _T_283; // @[Mux.scala 98:16]
  wire [1:0] _T_285 = _T_101 ? 2'h1 : _T_284; // @[Mux.scala 98:16]
  wire [1:0] _T_286 = _T_99 ? 2'h1 : _T_285; // @[Mux.scala 98:16]
  wire [1:0] _T_287 = _T_97 ? 2'h1 : _T_286; // @[Mux.scala 98:16]
  wire [1:0] _T_288 = _T_95 ? 2'h1 : _T_287; // @[Mux.scala 98:16]
  wire [1:0] _T_289 = _T_93 ? 2'h1 : _T_288; // @[Mux.scala 98:16]
  wire [1:0] _T_290 = _T_91 ? 2'h1 : _T_289; // @[Mux.scala 98:16]
  wire [1:0] _T_291 = _T_89 ? 2'h1 : _T_290; // @[Mux.scala 98:16]
  wire [1:0] _T_292 = _T_87 ? 2'h0 : _T_291; // @[Mux.scala 98:16]
  wire [1:0] _T_293 = _T_85 ? 2'h1 : _T_292; // @[Mux.scala 98:16]
  wire [1:0] _T_294 = _T_83 ? 2'h0 : _T_293; // @[Mux.scala 98:16]
  wire [1:0] _T_295 = _T_81 ? 2'h0 : _T_294; // @[Mux.scala 98:16]
  wire [1:0] _T_296 = _T_79 ? 2'h1 : _T_295; // @[Mux.scala 98:16]
  wire [1:0] _T_297 = _T_77 ? 2'h0 : _T_296; // @[Mux.scala 98:16]
  wire [1:0] _T_298 = _T_75 ? 2'h1 : _T_297; // @[Mux.scala 98:16]
  wire [1:0] _T_299 = _T_73 ? 2'h0 : _T_298; // @[Mux.scala 98:16]
  wire [1:0] _T_300 = _T_71 ? 2'h0 : _T_299; // @[Mux.scala 98:16]
  wire [1:0] _T_301 = _T_69 ? 2'h1 : _T_300; // @[Mux.scala 98:16]
  wire [1:0] _T_302 = _T_67 ? 2'h0 : _T_301; // @[Mux.scala 98:16]
  wire [1:0] _T_303 = _T_65 ? 2'h1 : _T_302; // @[Mux.scala 98:16]
  wire [1:0] _T_304 = _T_63 ? 2'h0 : _T_303; // @[Mux.scala 98:16]
  wire [1:0] _T_305 = _T_61 ? 2'h0 : _T_304; // @[Mux.scala 98:16]
  wire [1:0] _T_306 = _T_59 ? 2'h1 : _T_305; // @[Mux.scala 98:16]
  wire [1:0] _T_307 = _T_57 ? 2'h0 : _T_306; // @[Mux.scala 98:16]
  wire [1:0] _T_308 = _T_55 ? 2'h1 : _T_307; // @[Mux.scala 98:16]
  wire [1:0] _T_309 = _T_53 ? 2'h0 : _T_308; // @[Mux.scala 98:16]
  wire [1:0] _T_310 = _T_51 ? 2'h0 : _T_309; // @[Mux.scala 98:16]
  wire [1:0] _T_311 = _T_49 ? 2'h1 : _T_310; // @[Mux.scala 98:16]
  wire [1:0] _T_312 = _T_47 ? 2'h1 : _T_311; // @[Mux.scala 98:16]
  wire [1:0] _T_313 = _T_45 ? 2'h1 : _T_312; // @[Mux.scala 98:16]
  wire [1:0] _T_314 = _T_43 ? 2'h0 : _T_313; // @[Mux.scala 98:16]
  wire [1:0] _T_315 = _T_41 ? 2'h0 : _T_314; // @[Mux.scala 98:16]
  wire [1:0] _T_316 = _T_39 ? 2'h0 : _T_315; // @[Mux.scala 98:16]
  wire [1:0] _T_317 = _T_37 ? 2'h0 : _T_316; // @[Mux.scala 98:16]
  wire [1:0] _T_318 = _T_35 ? 2'h0 : _T_317; // @[Mux.scala 98:16]
  wire [1:0] _T_319 = _T_33 ? 2'h1 : _T_318; // @[Mux.scala 98:16]
  wire [1:0] _T_320 = _T_31 ? 2'h0 : _T_319; // @[Mux.scala 98:16]
  wire [1:0] _T_321 = _T_29 ? 2'h0 : _T_320; // @[Mux.scala 98:16]
  wire [1:0] _T_322 = _T_27 ? 2'h0 : _T_321; // @[Mux.scala 98:16]
  wire [1:0] _T_323 = _T_25 ? 2'h0 : _T_322; // @[Mux.scala 98:16]
  wire [1:0] _T_324 = _T_23 ? 2'h1 : _T_323; // @[Mux.scala 98:16]
  wire [1:0] _T_325 = _T_21 ? 2'h0 : _T_324; // @[Mux.scala 98:16]
  wire [1:0] _T_326 = _T_19 ? 2'h0 : _T_325; // @[Mux.scala 98:16]
  wire [1:0] _T_327 = _T_17 ? 2'h0 : _T_326; // @[Mux.scala 98:16]
  wire [1:0] _T_328 = _T_15 ? 2'h1 : _T_327; // @[Mux.scala 98:16]
  wire [1:0] _T_329 = _T_13 ? 2'h0 : _T_328; // @[Mux.scala 98:16]
  wire [1:0] _T_330 = _T_11 ? 2'h1 : _T_329; // @[Mux.scala 98:16]
  wire [1:0] _T_331 = _T_9 ? 2'h0 : _T_330; // @[Mux.scala 98:16]
  wire [1:0] _T_332 = _T_7 ? 2'h0 : _T_331; // @[Mux.scala 98:16]
  wire [1:0] _T_333 = _T_5 ? 2'h1 : _T_332; // @[Mux.scala 98:16]
  wire [1:0] _T_334 = _T_3 ? 2'h1 : _T_333; // @[Mux.scala 98:16]
  assign io_AluSrc1 = {{1'd0}, _T_279}; // @[ALUSrcGen.scala 91:14]
  assign io_AluSrc2 = _T_1 ? 2'h0 : _T_334; // @[ALUSrcGen.scala 92:14]
endmodule
module memWriteMGen(
  input  [31:0] io_inst,
  output        io_memWriteM
);
  wire [31:0] _T = io_inst & 32'h707f; // @[memWriteMGen.scala 20:49]
  wire  _T_1 = 32'h3023 == _T; // @[memWriteMGen.scala 20:49]
  wire  _T_3 = 32'h2023 == _T; // @[memWriteMGen.scala 20:49]
  wire  _T_5 = 32'h23 == _T; // @[memWriteMGen.scala 20:49]
  wire  _T_7 = 32'h1023 == _T; // @[memWriteMGen.scala 20:49]
  wire  _T_9 = _T_5 | _T_7; // @[Mux.scala 98:16]
  wire  _T_10 = _T_3 | _T_9; // @[Mux.scala 98:16]
  assign io_memWriteM = _T_1 | _T_10; // @[memWriteMGen.scala 26:16]
endmodule
module memWriteMaskGen(
  input  [31:0] io_inst,
  output [7:0]  io_mask
);
  wire  _T_1 = 3'h0 == io_inst[14:12]; // @[Mux.scala 80:60]
  wire [7:0] _T_2 = _T_1 ? 8'h1 : 8'h0; // @[Mux.scala 80:57]
  wire  _T_3 = 3'h1 == io_inst[14:12]; // @[Mux.scala 80:60]
  wire [7:0] _T_4 = _T_3 ? 8'h3 : _T_2; // @[Mux.scala 80:57]
  wire  _T_5 = 3'h2 == io_inst[14:12]; // @[Mux.scala 80:60]
  wire [7:0] _T_6 = _T_5 ? 8'hf : _T_4; // @[Mux.scala 80:57]
  wire  _T_7 = 3'h3 == io_inst[14:12]; // @[Mux.scala 80:60]
  assign io_mask = _T_7 ? 8'hff : _T_6; // @[memWriteMaskGen.scala 20:11]
endmodule
module memReadNumGen(
  input  [31:0] io_inst,
  output [2:0]  io_memReadNum
);
  assign io_memReadNum = io_inst[14:12]; // @[memReadNumGen.scala 23:17]
endmodule
module dnpcSrcGen(
  input  [31:0] io_inst,
  output        io_dnpcSrc
);
  wire [31:0] _T = io_inst & 32'h707f; // @[npcSrcGen.scala 26:49]
  wire  _T_1 = 32'h6063 == _T; // @[npcSrcGen.scala 26:49]
  wire  _T_3 = 32'h5063 == _T; // @[npcSrcGen.scala 26:49]
  wire  _T_5 = 32'h1063 == _T; // @[npcSrcGen.scala 26:49]
  wire  _T_7 = 32'h4063 == _T; // @[npcSrcGen.scala 26:49]
  wire  _T_9 = 32'h63 == _T; // @[npcSrcGen.scala 26:49]
  wire  _T_11 = 32'h7063 == _T; // @[npcSrcGen.scala 26:49]
  wire [31:0] _T_12 = io_inst & 32'h7f; // @[npcSrcGen.scala 31:31]
  wire  _T_13 = 32'h6f == _T_12; // @[npcSrcGen.scala 31:31]
  wire  _T_18 = _T_11 | _T_13; // @[Mux.scala 98:16]
  wire  _T_19 = _T_9 | _T_18; // @[Mux.scala 98:16]
  wire  _T_20 = _T_7 | _T_19; // @[Mux.scala 98:16]
  wire  _T_21 = _T_5 | _T_20; // @[Mux.scala 98:16]
  wire  _T_22 = _T_3 | _T_21; // @[Mux.scala 98:16]
  assign io_dnpcSrc = _T_1 | _T_22; // @[npcSrcGen.scala 34:14]
endmodule
module jumpGen(
  input  [31:0] io_inst,
  output        io_jump
);
  wire [31:0] _T = io_inst & 32'h7f; // @[npcSrcGen.scala 47:14]
  wire  _T_1 = 32'h6f == _T; // @[npcSrcGen.scala 47:14]
  wire [31:0] _T_2 = io_inst & 32'h707f; // @[npcSrcGen.scala 48:14]
  wire  _T_3 = 32'h67 == _T_2; // @[npcSrcGen.scala 48:14]
  assign io_jump = _T_1 | _T_3; // @[npcSrcGen.scala 51:11]
endmodule
module branchGen(
  input  [31:0] io_inst,
  output        io_branch
);
  wire [31:0] _T = io_inst & 32'h707f; // @[npcSrcGen.scala 67:47]
  wire  _T_1 = 32'h6063 == _T; // @[npcSrcGen.scala 67:47]
  wire  _T_3 = 32'h5063 == _T; // @[npcSrcGen.scala 67:47]
  wire  _T_5 = 32'h1063 == _T; // @[npcSrcGen.scala 67:47]
  wire  _T_7 = 32'h4063 == _T; // @[npcSrcGen.scala 67:47]
  wire  _T_9 = 32'h63 == _T; // @[npcSrcGen.scala 67:47]
  wire  _T_11 = 32'h7063 == _T; // @[npcSrcGen.scala 67:47]
  wire  _T_13 = _T_9 | _T_11; // @[Mux.scala 98:16]
  wire  _T_14 = _T_7 | _T_13; // @[Mux.scala 98:16]
  wire  _T_15 = _T_5 | _T_14; // @[Mux.scala 98:16]
  wire  _T_16 = _T_3 | _T_15; // @[Mux.scala 98:16]
  assign io_branch = _T_1 | _T_16; // @[npcSrcGen.scala 73:13]
endmodule
module regEnGen(
  input  [31:0] io_inst,
  output        io_regEn
);
  wire [31:0] _T = io_inst & 32'hfe00707f; // @[regEnGen.scala 35:45]
  wire  _T_1 = 32'h4033 == _T; // @[regEnGen.scala 35:45]
  wire [31:0] _T_2 = io_inst & 32'h707f; // @[regEnGen.scala 36:45]
  wire  _T_3 = 32'h3023 == _T_2; // @[regEnGen.scala 36:45]
  wire [31:0] _T_4 = io_inst & 32'hfc00707f; // @[regEnGen.scala 33:45]
  wire  _T_5 = 32'h1013 == _T_4; // @[regEnGen.scala 33:45]
  wire  _T_7 = 32'h503b == _T; // @[regEnGen.scala 35:45]
  wire  _T_9 = 32'h6063 == _T_2; // @[regEnGen.scala 37:45]
  wire  _T_11 = 32'h1003 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_13 = 32'h2004033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_15 = 32'h4013 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_17 = 32'h2006033 == _T; // @[regEnGen.scala 35:45]
  wire [31:0] _T_18 = io_inst & 32'h7f; // @[regEnGen.scala 34:45]
  wire  _T_19 = 32'h6f == _T_18; // @[regEnGen.scala 34:45]
  wire  _T_21 = 32'h200403b == _T; // @[regEnGen.scala 35:45]
  wire  _T_23 = 32'h3033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_25 = 32'h6013 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_27 = 32'h5033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_29 = 32'h5063 == _T_2; // @[regEnGen.scala 37:45]
  wire  _T_31 = 32'h6033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_33 = 32'h4000503b == _T; // @[regEnGen.scala 35:45]
  wire  _T_35 = 32'h7013 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_37 = 32'h33 == _T; // @[regEnGen.scala 35:45]
  wire  _T_39 = 32'h103b == _T; // @[regEnGen.scala 35:45]
  wire  _T_41 = 32'h2000033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_43 = 32'h2005033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_45 = 32'h2033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_47 = 32'h4003 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_49 = 32'h3 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_51 = 32'h2023 == _T_2; // @[regEnGen.scala 36:45]
  wire  _T_53 = 32'h200703b == _T; // @[regEnGen.scala 35:45]
  wire  _T_55 = 32'h1063 == _T_2; // @[regEnGen.scala 37:45]
  wire  _T_57 = 32'h1b == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_59 = 32'h17 == _T_18; // @[regEnGen.scala 32:45]
  wire  _T_61 = 32'h4063 == _T_2; // @[regEnGen.scala 37:45]
  wire  _T_63 = 32'h40005013 == _T_4; // @[regEnGen.scala 33:45]
  wire  _T_65 = 32'h200603b == _T; // @[regEnGen.scala 35:45]
  wire  _T_67 = 32'h63 == _T_2; // @[regEnGen.scala 37:45]
  wire  _T_69 = 32'h3003 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_71 = 32'h3b == _T; // @[regEnGen.scala 35:45]
  wire  _T_73 = 32'h4000501b == _T; // @[regEnGen.scala 33:45]
  wire  _T_75 = 32'h7033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_77 = 32'h200003b == _T; // @[regEnGen.scala 35:45]
  wire  _T_79 = 32'h67 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_81 = 32'h2007033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_83 = 32'h5013 == _T_4; // @[regEnGen.scala 33:45]
  wire  _T_85 = 32'h4000003b == _T; // @[regEnGen.scala 35:45]
  wire  _T_87 = 32'h200503b == _T; // @[regEnGen.scala 35:45]
  wire  _T_89 = 32'h23 == _T_2; // @[regEnGen.scala 36:45]
  wire  _T_91 = 32'h37 == _T_18; // @[regEnGen.scala 32:45]
  wire  _T_93 = 32'h40000033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_95 = 32'h501b == _T; // @[regEnGen.scala 33:45]
  wire  _T_97 = 32'h5003 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_99 = 32'h6003 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_101 = 32'h2003 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_103 = 32'h101b == _T; // @[regEnGen.scala 33:45]
  wire  _T_105 = 32'h1023 == _T_2; // @[regEnGen.scala 36:45]
  wire  _T_107 = 32'h13 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_109 = 32'h7063 == _T_2; // @[regEnGen.scala 37:45]
  wire  _T_111 = 32'h1033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_113 = 32'h3013 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_115 = _T_111 | _T_113; // @[Mux.scala 98:16]
  wire  _T_116 = _T_109 ? 1'h0 : _T_115; // @[Mux.scala 98:16]
  wire  _T_117 = _T_107 | _T_116; // @[Mux.scala 98:16]
  wire  _T_118 = _T_105 ? 1'h0 : _T_117; // @[Mux.scala 98:16]
  wire  _T_119 = _T_103 | _T_118; // @[Mux.scala 98:16]
  wire  _T_120 = _T_101 | _T_119; // @[Mux.scala 98:16]
  wire  _T_121 = _T_99 | _T_120; // @[Mux.scala 98:16]
  wire  _T_122 = _T_97 | _T_121; // @[Mux.scala 98:16]
  wire  _T_123 = _T_95 | _T_122; // @[Mux.scala 98:16]
  wire  _T_124 = _T_93 | _T_123; // @[Mux.scala 98:16]
  wire  _T_125 = _T_91 | _T_124; // @[Mux.scala 98:16]
  wire  _T_126 = _T_89 ? 1'h0 : _T_125; // @[Mux.scala 98:16]
  wire  _T_127 = _T_87 | _T_126; // @[Mux.scala 98:16]
  wire  _T_128 = _T_85 | _T_127; // @[Mux.scala 98:16]
  wire  _T_129 = _T_83 | _T_128; // @[Mux.scala 98:16]
  wire  _T_130 = _T_81 | _T_129; // @[Mux.scala 98:16]
  wire  _T_131 = _T_79 | _T_130; // @[Mux.scala 98:16]
  wire  _T_132 = _T_77 | _T_131; // @[Mux.scala 98:16]
  wire  _T_133 = _T_75 | _T_132; // @[Mux.scala 98:16]
  wire  _T_134 = _T_73 | _T_133; // @[Mux.scala 98:16]
  wire  _T_135 = _T_71 | _T_134; // @[Mux.scala 98:16]
  wire  _T_136 = _T_69 | _T_135; // @[Mux.scala 98:16]
  wire  _T_137 = _T_67 ? 1'h0 : _T_136; // @[Mux.scala 98:16]
  wire  _T_138 = _T_65 | _T_137; // @[Mux.scala 98:16]
  wire  _T_139 = _T_63 | _T_138; // @[Mux.scala 98:16]
  wire  _T_140 = _T_61 ? 1'h0 : _T_139; // @[Mux.scala 98:16]
  wire  _T_141 = _T_59 | _T_140; // @[Mux.scala 98:16]
  wire  _T_142 = _T_57 | _T_141; // @[Mux.scala 98:16]
  wire  _T_143 = _T_55 ? 1'h0 : _T_142; // @[Mux.scala 98:16]
  wire  _T_144 = _T_53 | _T_143; // @[Mux.scala 98:16]
  wire  _T_145 = _T_51 ? 1'h0 : _T_144; // @[Mux.scala 98:16]
  wire  _T_146 = _T_49 | _T_145; // @[Mux.scala 98:16]
  wire  _T_147 = _T_47 | _T_146; // @[Mux.scala 98:16]
  wire  _T_148 = _T_45 | _T_147; // @[Mux.scala 98:16]
  wire  _T_149 = _T_43 | _T_148; // @[Mux.scala 98:16]
  wire  _T_150 = _T_41 | _T_149; // @[Mux.scala 98:16]
  wire  _T_151 = _T_39 | _T_150; // @[Mux.scala 98:16]
  wire  _T_152 = _T_37 | _T_151; // @[Mux.scala 98:16]
  wire  _T_153 = _T_35 | _T_152; // @[Mux.scala 98:16]
  wire  _T_154 = _T_33 | _T_153; // @[Mux.scala 98:16]
  wire  _T_155 = _T_31 | _T_154; // @[Mux.scala 98:16]
  wire  _T_156 = _T_29 ? 1'h0 : _T_155; // @[Mux.scala 98:16]
  wire  _T_157 = _T_27 | _T_156; // @[Mux.scala 98:16]
  wire  _T_158 = _T_25 | _T_157; // @[Mux.scala 98:16]
  wire  _T_159 = _T_23 | _T_158; // @[Mux.scala 98:16]
  wire  _T_160 = _T_21 | _T_159; // @[Mux.scala 98:16]
  wire  _T_161 = _T_19 | _T_160; // @[Mux.scala 98:16]
  wire  _T_162 = _T_17 | _T_161; // @[Mux.scala 98:16]
  wire  _T_163 = _T_15 | _T_162; // @[Mux.scala 98:16]
  wire  _T_164 = _T_13 | _T_163; // @[Mux.scala 98:16]
  wire  _T_165 = _T_11 | _T_164; // @[Mux.scala 98:16]
  wire  _T_166 = _T_9 ? 1'h0 : _T_165; // @[Mux.scala 98:16]
  wire  _T_167 = _T_7 | _T_166; // @[Mux.scala 98:16]
  wire  _T_168 = _T_5 | _T_167; // @[Mux.scala 98:16]
  wire  _T_169 = _T_3 ? 1'h0 : _T_168; // @[Mux.scala 98:16]
  assign io_regEn = _T_1 | _T_169; // @[regEnGen.scala 43:12]
endmodule
module ResultSrcGen(
  input  [31:0] io_inst,
  output [1:0]  io_ResultSrc
);
  wire [31:0] _T = io_inst & 32'hfe00707f; // @[ResultSrcGen.scala 40:44]
  wire  _T_1 = 32'h4033 == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_3 = 32'h503b == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_5 = 32'h2004033 == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_7 = 32'h2006033 == _T; // @[ResultSrcGen.scala 40:44]
  wire [31:0] _T_8 = io_inst & 32'h7f; // @[ResultSrcGen.scala 39:44]
  wire  _T_9 = 32'h6f == _T_8; // @[ResultSrcGen.scala 39:44]
  wire  _T_11 = 32'h200403b == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_13 = 32'h3033 == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_15 = 32'h5033 == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_17 = 32'h6033 == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_19 = 32'h4000503b == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_21 = 32'h33 == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_23 = 32'h103b == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_25 = 32'h2000033 == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_27 = 32'h2005033 == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_29 = 32'h2033 == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_31 = 32'h200703b == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_33 = 32'h17 == _T_8; // @[ResultSrcGen.scala 38:44]
  wire  _T_35 = 32'h200603b == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_37 = 32'h3b == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_39 = 32'h7033 == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_41 = 32'h200003b == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_43 = 32'h2007033 == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_45 = 32'h4000003b == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_47 = 32'h200503b == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_49 = 32'h37 == _T_8; // @[ResultSrcGen.scala 38:44]
  wire  _T_51 = 32'h40000033 == _T; // @[ResultSrcGen.scala 40:44]
  wire  _T_53 = 32'h1033 == _T; // @[ResultSrcGen.scala 40:44]
  wire [31:0] _T_54 = io_inst & 32'h707f; // @[ResultSrcGen.scala 45:26]
  wire  _T_55 = 32'h13 == _T_54; // @[ResultSrcGen.scala 45:26]
  wire  _T_57 = 32'h67 == _T_54; // @[ResultSrcGen.scala 46:26]
  wire  _T_61 = 32'h3003 == _T_54; // @[ResultSrcGen.scala 48:26]
  wire  _T_63 = 32'h4003 == _T_54; // @[ResultSrcGen.scala 49:26]
  wire  _T_65 = 32'h3013 == _T_54; // @[ResultSrcGen.scala 50:26]
  wire  _T_67 = 32'h501b == _T; // @[ResultSrcGen.scala 51:26]
  wire [31:0] _T_68 = io_inst & 32'hfc00707f; // @[ResultSrcGen.scala 52:26]
  wire  _T_69 = 32'h1013 == _T_68; // @[ResultSrcGen.scala 52:26]
  wire  _T_71 = 32'h7013 == _T_54; // @[ResultSrcGen.scala 53:26]
  wire  _T_73 = 32'h4013 == _T_54; // @[ResultSrcGen.scala 54:26]
  wire  _T_75 = 32'h1b == _T_54; // @[ResultSrcGen.scala 55:26]
  wire  _T_77 = 32'h5013 == _T_68; // @[ResultSrcGen.scala 56:26]
  wire  _T_79 = 32'h101b == _T; // @[ResultSrcGen.scala 57:26]
  wire  _T_81 = 32'h4000501b == _T; // @[ResultSrcGen.scala 58:26]
  wire  _T_83 = 32'h40005013 == _T_68; // @[ResultSrcGen.scala 59:26]
  wire  _T_85 = 32'h6013 == _T_54; // @[ResultSrcGen.scala 60:26]
  wire  _T_87 = 32'h1003 == _T_54; // @[ResultSrcGen.scala 61:26]
  wire  _T_89 = 32'h2003 == _T_54; // @[ResultSrcGen.scala 62:26]
  wire  _T_91 = 32'h5003 == _T_54; // @[ResultSrcGen.scala 63:26]
  wire  _T_93 = 32'h6003 == _T_54; // @[ResultSrcGen.scala 64:26]
  wire  _T_95 = 32'h3 == _T_54; // @[ResultSrcGen.scala 65:26]
  wire [1:0] _T_102 = _T_95 ? 2'h2 : 2'h0; // @[Mux.scala 98:16]
  wire [1:0] _T_103 = _T_93 ? 2'h2 : _T_102; // @[Mux.scala 98:16]
  wire [1:0] _T_104 = _T_91 ? 2'h2 : _T_103; // @[Mux.scala 98:16]
  wire [1:0] _T_105 = _T_89 ? 2'h2 : _T_104; // @[Mux.scala 98:16]
  wire [1:0] _T_106 = _T_87 ? 2'h2 : _T_105; // @[Mux.scala 98:16]
  wire [1:0] _T_107 = _T_85 ? 2'h0 : _T_106; // @[Mux.scala 98:16]
  wire [1:0] _T_108 = _T_83 ? 2'h0 : _T_107; // @[Mux.scala 98:16]
  wire [1:0] _T_109 = _T_81 ? 2'h0 : _T_108; // @[Mux.scala 98:16]
  wire [1:0] _T_110 = _T_79 ? 2'h0 : _T_109; // @[Mux.scala 98:16]
  wire [1:0] _T_111 = _T_77 ? 2'h0 : _T_110; // @[Mux.scala 98:16]
  wire [1:0] _T_112 = _T_75 ? 2'h0 : _T_111; // @[Mux.scala 98:16]
  wire [1:0] _T_113 = _T_73 ? 2'h0 : _T_112; // @[Mux.scala 98:16]
  wire [1:0] _T_114 = _T_71 ? 2'h0 : _T_113; // @[Mux.scala 98:16]
  wire [1:0] _T_115 = _T_69 ? 2'h0 : _T_114; // @[Mux.scala 98:16]
  wire [1:0] _T_116 = _T_67 ? 2'h0 : _T_115; // @[Mux.scala 98:16]
  wire [1:0] _T_117 = _T_65 ? 2'h0 : _T_116; // @[Mux.scala 98:16]
  wire [1:0] _T_118 = _T_63 ? 2'h2 : _T_117; // @[Mux.scala 98:16]
  wire [1:0] _T_119 = _T_61 ? 2'h2 : _T_118; // @[Mux.scala 98:16]
  wire [1:0] _T_120 = _T_57 ? 2'h1 : _T_119; // @[Mux.scala 98:16]
  wire [1:0] _T_121 = _T_57 ? 2'h1 : _T_120; // @[Mux.scala 98:16]
  wire [1:0] _T_122 = _T_55 ? 2'h0 : _T_121; // @[Mux.scala 98:16]
  wire [1:0] _T_123 = _T_53 ? 2'h0 : _T_122; // @[Mux.scala 98:16]
  wire [1:0] _T_124 = _T_51 ? 2'h0 : _T_123; // @[Mux.scala 98:16]
  wire [1:0] _T_125 = _T_49 ? 2'h0 : _T_124; // @[Mux.scala 98:16]
  wire [1:0] _T_126 = _T_47 ? 2'h0 : _T_125; // @[Mux.scala 98:16]
  wire [1:0] _T_127 = _T_45 ? 2'h0 : _T_126; // @[Mux.scala 98:16]
  wire [1:0] _T_128 = _T_43 ? 2'h0 : _T_127; // @[Mux.scala 98:16]
  wire [1:0] _T_129 = _T_41 ? 2'h0 : _T_128; // @[Mux.scala 98:16]
  wire [1:0] _T_130 = _T_39 ? 2'h0 : _T_129; // @[Mux.scala 98:16]
  wire [1:0] _T_131 = _T_37 ? 2'h0 : _T_130; // @[Mux.scala 98:16]
  wire [1:0] _T_132 = _T_35 ? 2'h0 : _T_131; // @[Mux.scala 98:16]
  wire [1:0] _T_133 = _T_33 ? 2'h0 : _T_132; // @[Mux.scala 98:16]
  wire [1:0] _T_134 = _T_31 ? 2'h0 : _T_133; // @[Mux.scala 98:16]
  wire [1:0] _T_135 = _T_29 ? 2'h0 : _T_134; // @[Mux.scala 98:16]
  wire [1:0] _T_136 = _T_27 ? 2'h0 : _T_135; // @[Mux.scala 98:16]
  wire [1:0] _T_137 = _T_25 ? 2'h0 : _T_136; // @[Mux.scala 98:16]
  wire [1:0] _T_138 = _T_23 ? 2'h0 : _T_137; // @[Mux.scala 98:16]
  wire [1:0] _T_139 = _T_21 ? 2'h0 : _T_138; // @[Mux.scala 98:16]
  wire [1:0] _T_140 = _T_19 ? 2'h0 : _T_139; // @[Mux.scala 98:16]
  wire [1:0] _T_141 = _T_17 ? 2'h0 : _T_140; // @[Mux.scala 98:16]
  wire [1:0] _T_142 = _T_15 ? 2'h0 : _T_141; // @[Mux.scala 98:16]
  wire [1:0] _T_143 = _T_13 ? 2'h0 : _T_142; // @[Mux.scala 98:16]
  wire [1:0] _T_144 = _T_11 ? 2'h0 : _T_143; // @[Mux.scala 98:16]
  wire [1:0] _T_145 = _T_9 ? 2'h1 : _T_144; // @[Mux.scala 98:16]
  wire [1:0] _T_146 = _T_7 ? 2'h0 : _T_145; // @[Mux.scala 98:16]
  wire [1:0] _T_147 = _T_5 ? 2'h0 : _T_146; // @[Mux.scala 98:16]
  wire [1:0] _T_148 = _T_3 ? 2'h0 : _T_147; // @[Mux.scala 98:16]
  assign io_ResultSrc = _T_1 ? 2'h0 : _T_148; // @[ResultSrcGen.scala 69:16]
endmodule
module CtrlUnit(
  input  [31:0] io_inst,
  output [1:0]  io_CtrlS_AluSrc1,
  output [1:0]  io_CtrlS_AluSrc2,
  output [4:0]  io_CtrlS_ALUCtrl,
  output        io_CtrlS_memWriteM,
  output [7:0]  io_CtrlS_memWriteMask,
  output [2:0]  io_CtrlS_memReadNum,
  output        io_CtrlS_dnpcSrc,
  output        io_CtrlS_jump,
  output        io_CtrlS_branch,
  output        io_CtrlS_regEn,
  output [1:0]  io_CtrlS_ResultSrc,
  output        io_CtrlS_fencei
);
  wire [31:0] ALUCtrl_ins_io_inst; // @[CtrlUnit.scala 33:26]
  wire [4:0] ALUCtrl_ins_io_ALUCtrl; // @[CtrlUnit.scala 33:26]
  wire [31:0] ALUSrcGen_ins_io_inst; // @[CtrlUnit.scala 37:29]
  wire [1:0] ALUSrcGen_ins_io_AluSrc1; // @[CtrlUnit.scala 37:29]
  wire [1:0] ALUSrcGen_ins_io_AluSrc2; // @[CtrlUnit.scala 37:29]
  wire [31:0] memWriteMGen_ins_io_inst; // @[CtrlUnit.scala 42:32]
  wire  memWriteMGen_ins_io_memWriteM; // @[CtrlUnit.scala 42:32]
  wire [31:0] memWriteMaskGen_ins_io_inst; // @[CtrlUnit.scala 46:35]
  wire [7:0] memWriteMaskGen_ins_io_mask; // @[CtrlUnit.scala 46:35]
  wire [31:0] memReadNumGen_ins_io_inst; // @[CtrlUnit.scala 50:33]
  wire [2:0] memReadNumGen_ins_io_memReadNum; // @[CtrlUnit.scala 50:33]
  wire [31:0] dnpcSrcGen_ins_io_inst; // @[CtrlUnit.scala 54:32]
  wire  dnpcSrcGen_ins_io_dnpcSrc; // @[CtrlUnit.scala 54:32]
  wire [31:0] jumpGen_ins_io_inst; // @[CtrlUnit.scala 58:27]
  wire  jumpGen_ins_io_jump; // @[CtrlUnit.scala 58:27]
  wire [31:0] branchGen_ins_io_inst; // @[CtrlUnit.scala 62:29]
  wire  branchGen_ins_io_branch; // @[CtrlUnit.scala 62:29]
  wire [31:0] regEnGen_ins_io_inst; // @[CtrlUnit.scala 67:28]
  wire  regEnGen_ins_io_regEn; // @[CtrlUnit.scala 67:28]
  wire [31:0] ResultSrcGen_ins_io_inst; // @[CtrlUnit.scala 71:32]
  wire [1:0] ResultSrcGen_ins_io_ResultSrc; // @[CtrlUnit.scala 71:32]
  wire [31:0] _T = io_inst & 32'h707f; // @[CtrlUnit.scala 75:30]
  ALUCtrl ALUCtrl_ins ( // @[CtrlUnit.scala 33:26]
    .io_inst(ALUCtrl_ins_io_inst),
    .io_ALUCtrl(ALUCtrl_ins_io_ALUCtrl)
  );
  ALUSrcGen ALUSrcGen_ins ( // @[CtrlUnit.scala 37:29]
    .io_inst(ALUSrcGen_ins_io_inst),
    .io_AluSrc1(ALUSrcGen_ins_io_AluSrc1),
    .io_AluSrc2(ALUSrcGen_ins_io_AluSrc2)
  );
  memWriteMGen memWriteMGen_ins ( // @[CtrlUnit.scala 42:32]
    .io_inst(memWriteMGen_ins_io_inst),
    .io_memWriteM(memWriteMGen_ins_io_memWriteM)
  );
  memWriteMaskGen memWriteMaskGen_ins ( // @[CtrlUnit.scala 46:35]
    .io_inst(memWriteMaskGen_ins_io_inst),
    .io_mask(memWriteMaskGen_ins_io_mask)
  );
  memReadNumGen memReadNumGen_ins ( // @[CtrlUnit.scala 50:33]
    .io_inst(memReadNumGen_ins_io_inst),
    .io_memReadNum(memReadNumGen_ins_io_memReadNum)
  );
  dnpcSrcGen dnpcSrcGen_ins ( // @[CtrlUnit.scala 54:32]
    .io_inst(dnpcSrcGen_ins_io_inst),
    .io_dnpcSrc(dnpcSrcGen_ins_io_dnpcSrc)
  );
  jumpGen jumpGen_ins ( // @[CtrlUnit.scala 58:27]
    .io_inst(jumpGen_ins_io_inst),
    .io_jump(jumpGen_ins_io_jump)
  );
  branchGen branchGen_ins ( // @[CtrlUnit.scala 62:29]
    .io_inst(branchGen_ins_io_inst),
    .io_branch(branchGen_ins_io_branch)
  );
  regEnGen regEnGen_ins ( // @[CtrlUnit.scala 67:28]
    .io_inst(regEnGen_ins_io_inst),
    .io_regEn(regEnGen_ins_io_regEn)
  );
  ResultSrcGen ResultSrcGen_ins ( // @[CtrlUnit.scala 71:32]
    .io_inst(ResultSrcGen_ins_io_inst),
    .io_ResultSrc(ResultSrcGen_ins_io_ResultSrc)
  );
  assign io_CtrlS_AluSrc1 = ALUSrcGen_ins_io_AluSrc1; // @[CtrlUnit.scala 39:20]
  assign io_CtrlS_AluSrc2 = ALUSrcGen_ins_io_AluSrc2; // @[CtrlUnit.scala 40:20]
  assign io_CtrlS_ALUCtrl = ALUCtrl_ins_io_ALUCtrl; // @[CtrlUnit.scala 35:20]
  assign io_CtrlS_memWriteM = memWriteMGen_ins_io_memWriteM; // @[CtrlUnit.scala 44:22]
  assign io_CtrlS_memWriteMask = memWriteMaskGen_ins_io_mask; // @[CtrlUnit.scala 48:25]
  assign io_CtrlS_memReadNum = memReadNumGen_ins_io_memReadNum; // @[CtrlUnit.scala 52:23]
  assign io_CtrlS_dnpcSrc = dnpcSrcGen_ins_io_dnpcSrc; // @[CtrlUnit.scala 56:20]
  assign io_CtrlS_jump = jumpGen_ins_io_jump; // @[CtrlUnit.scala 60:17]
  assign io_CtrlS_branch = branchGen_ins_io_branch; // @[CtrlUnit.scala 64:19]
  assign io_CtrlS_regEn = regEnGen_ins_io_regEn; // @[CtrlUnit.scala 69:18]
  assign io_CtrlS_ResultSrc = ResultSrcGen_ins_io_ResultSrc; // @[CtrlUnit.scala 73:22]
  assign io_CtrlS_fencei = 32'h100f == _T; // @[CtrlUnit.scala 75:19]
  assign ALUCtrl_ins_io_inst = io_inst; // @[CtrlUnit.scala 34:23]
  assign ALUSrcGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 38:25]
  assign memWriteMGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 43:28]
  assign memWriteMaskGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 47:31]
  assign memReadNumGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 51:29]
  assign dnpcSrcGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 55:26]
  assign jumpGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 59:23]
  assign branchGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 63:25]
  assign regEnGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 68:24]
  assign ResultSrcGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 72:28]
endmodule
module csrCtrl(
  input  [31:0] io_inst,
  output        io_CSRCtrlIf_csrrwen,
  output        io_CSRCtrlIf_csrswen,
  output        io_CSRCtrlIf_csrrsien,
  output        io_CSRCtrlIf_csrrcien,
  output        io_CSRCtrlIf_csrrcen,
  output        io_CSRCtrlIf_csrrwien,
  output        io_CSRCtrlIf_ecall,
  output        io_CSRCtrlIf_rfen,
  output        io_CSRCtrlIf_mepc2pc
);
  wire [31:0] _T_2 = io_inst & 32'h707f; // @[csrCtrl.scala 44:35]
  wire  _T_3 = 32'h1073 == _T_2; // @[csrCtrl.scala 44:35]
  wire  _T_5 = 32'h2073 == _T_2; // @[csrCtrl.scala 45:35]
  wire  _T_7 = 32'h6073 == _T_2; // @[csrCtrl.scala 46:36]
  wire  _T_9 = 32'h7073 == _T_2; // @[csrCtrl.scala 47:36]
  wire  _T_11 = 32'h3073 == _T_2; // @[csrCtrl.scala 48:35]
  wire  _T_18 = _T_3 | _T_5; // @[csrCtrl.scala 51:41]
  wire  _T_21 = _T_18 | _T_7; // @[csrCtrl.scala 51:61]
  wire  _T_24 = _T_21 | _T_9; // @[csrCtrl.scala 51:81]
  assign io_CSRCtrlIf_csrrwen = 32'h1073 == _T_2; // @[csrCtrl.scala 44:24]
  assign io_CSRCtrlIf_csrswen = 32'h2073 == _T_2; // @[csrCtrl.scala 45:24]
  assign io_CSRCtrlIf_csrrsien = 32'h6073 == _T_2; // @[csrCtrl.scala 46:25]
  assign io_CSRCtrlIf_csrrcien = 32'h7073 == _T_2; // @[csrCtrl.scala 47:25]
  assign io_CSRCtrlIf_csrrcen = 32'h3073 == _T_2; // @[csrCtrl.scala 48:24]
  assign io_CSRCtrlIf_csrrwien = 32'h5073 == _T_2; // @[csrCtrl.scala 49:25]
  assign io_CSRCtrlIf_ecall = 32'h73 == io_inst; // @[csrCtrl.scala 41:22]
  assign io_CSRCtrlIf_rfen = _T_24 | _T_11; // @[csrCtrl.scala 51:21]
  assign io_CSRCtrlIf_mepc2pc = 32'h30200073 == io_inst; // @[csrCtrl.scala 53:24]
endmodule
module riscv(
  input          clock,
  input          reset,
  output         io_instIO_valid,
  input          io_instIO_ready,
  input  [63:0]  io_instIO_data_read,
  output [31:0]  io_instIO_addr,
  output         io_dataIO_valid,
  input          io_dataIO_ready,
  input  [63:0]  io_dataIO_data_read,
  output [63:0]  io_dataIO_data_write,
  output         io_dataIO_wen,
  output [31:0]  io_dataIO_addr,
  output [1:0]   io_dataIO_rsize,
  output [7:0]   io_dataIO_mask,
  output         _T_99_0,
  input          intrTimeCnt_0,
  output         _T_100_0,
  output         startTimeCnt,
  output         block3_0,
  output [191:0] dmaCtrl,
  output         block2_0,
  input          blockDMA_0,
  output         fencei_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [287:0] _RAND_0;
  reg [447:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [191:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [95:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  ifu_clock; // @[riscv.scala 34:19]
  wire  ifu_reset; // @[riscv.scala 34:19]
  wire [31:0] ifu_io_instIn; // @[riscv.scala 34:19]
  wire [31:0] ifu_io_instOut; // @[riscv.scala 34:19]
  wire [31:0] ifu_io_pc; // @[riscv.scala 34:19]
  wire [31:0] ifu_io_snpc; // @[riscv.scala 34:19]
  wire [31:0] ifu_io_dnpc; // @[riscv.scala 34:19]
  wire  ifu_io_jump; // @[riscv.scala 34:19]
  wire  ifu_intrTimeCnt_0; // @[riscv.scala 34:19]
  wire  ifu_hazardPCBlock_0; // @[riscv.scala 34:19]
  wire  ifu_blockDMA_0; // @[riscv.scala 34:19]
  wire  ifu_block23_0; // @[riscv.scala 34:19]
  wire  ifu_block1_0; // @[riscv.scala 34:19]
  wire  idu_clock; // @[riscv.scala 35:19]
  wire  idu_reset; // @[riscv.scala 35:19]
  wire [31:0] idu_io_pc; // @[riscv.scala 35:19]
  wire [31:0] idu_io_inst; // @[riscv.scala 35:19]
  wire  idu_io_regEn; // @[riscv.scala 35:19]
  wire [63:0] idu_io_dataEx_imme; // @[riscv.scala 35:19]
  wire [63:0] idu_io_dataEx_dOut1; // @[riscv.scala 35:19]
  wire [63:0] idu_io_dataEx_dOut2; // @[riscv.scala 35:19]
  wire [63:0] idu_io_dataEx_dIn; // @[riscv.scala 35:19]
  wire [63:0] idu_io_dataEx_rdDout; // @[riscv.scala 35:19]
  wire [4:0] idu_io_rdOut; // @[riscv.scala 35:19]
  wire [4:0] idu_io_rdIn; // @[riscv.scala 35:19]
  wire [4:0] idu_io_rs1; // @[riscv.scala 35:19]
  wire [4:0] idu_io_rs2; // @[riscv.scala 35:19]
  wire [63:0] idu_io_dOutWB; // @[riscv.scala 35:19]
  wire  idu_blockDMA; // @[riscv.scala 35:19]
  wire  idu_block23; // @[riscv.scala 35:19]
  wire  idu_block1; // @[riscv.scala 35:19]
  wire  exu_clock; // @[riscv.scala 36:19]
  wire  exu_reset; // @[riscv.scala 36:19]
  wire [1:0] exu_io_AluSrc1; // @[riscv.scala 36:19]
  wire [1:0] exu_io_AluSrc2; // @[riscv.scala 36:19]
  wire [4:0] exu_io_ALUCtrl; // @[riscv.scala 36:19]
  wire  exu_io_dnpcSrc; // @[riscv.scala 36:19]
  wire [1:0] exu_io_ResultSrc; // @[riscv.scala 36:19]
  wire [2:0] exu_io_memReadNum; // @[riscv.scala 36:19]
  wire [63:0] exu_io_dataId_imme; // @[riscv.scala 36:19]
  wire [63:0] exu_io_dataId_dOut1; // @[riscv.scala 36:19]
  wire [63:0] exu_io_dataId_dOut2; // @[riscv.scala 36:19]
  wire [63:0] exu_io_dataId_dIn; // @[riscv.scala 36:19]
  wire [63:0] exu_io_dataId_rdDout; // @[riscv.scala 36:19]
  wire [63:0] exu_io_dataOut_ALUResOut; // @[riscv.scala 36:19]
  wire [63:0] exu_io_dataOut_wdata; // @[riscv.scala 36:19]
  wire [63:0] exu_io_dataOut_rdata; // @[riscv.scala 36:19]
  wire  exu_io_brTake; // @[riscv.scala 36:19]
  wire [31:0] exu_io_pc; // @[riscv.scala 36:19]
  wire [31:0] exu_io_snpc; // @[riscv.scala 36:19]
  wire [31:0] exu_io_dnpc; // @[riscv.scala 36:19]
  wire  exu_io_CSRCtrlIf_csrrwen; // @[riscv.scala 36:19]
  wire  exu_io_CSRCtrlIf_csrswen; // @[riscv.scala 36:19]
  wire  exu_io_CSRCtrlIf_csrrsien; // @[riscv.scala 36:19]
  wire  exu_io_CSRCtrlIf_csrrcien; // @[riscv.scala 36:19]
  wire  exu_io_CSRCtrlIf_csrrcen; // @[riscv.scala 36:19]
  wire  exu_io_CSRCtrlIf_csrrwien; // @[riscv.scala 36:19]
  wire  exu_io_CSRCtrlIf_ecall; // @[riscv.scala 36:19]
  wire  exu_io_CSRCtrlIf_rfen; // @[riscv.scala 36:19]
  wire  exu_io_CSRCtrlIf_mepc2pc; // @[riscv.scala 36:19]
  wire [4:0] exu_io_uimm; // @[riscv.scala 36:19]
  wire [63:0] exu_io_aluResIn; // @[riscv.scala 36:19]
  wire [1:0] exu_io_forwardA; // @[riscv.scala 36:19]
  wire [1:0] exu_io_forwardB; // @[riscv.scala 36:19]
  wire [1:0] exu_io_forwardC; // @[riscv.scala 36:19]
  wire [63:0] exu_io_aluRes1; // @[riscv.scala 36:19]
  wire [63:0] exu_io_aluRes3; // @[riscv.scala 36:19]
  wire  exu_intrTimeCnt_0; // @[riscv.scala 36:19]
  wire  exu_startTimeCnt; // @[riscv.scala 36:19]
  wire [191:0] exu_dmaCtrl_0; // @[riscv.scala 36:19]
  wire  exu_blockDMA; // @[riscv.scala 36:19]
  wire  exu_block23; // @[riscv.scala 36:19]
  wire  exu_block1; // @[riscv.scala 36:19]
  wire  hazardu_io_regEnEXMEM; // @[riscv.scala 37:23]
  wire [4:0] hazardu_io_rdEXMEM; // @[riscv.scala 37:23]
  wire [4:0] hazardu_io_rs1IDEX; // @[riscv.scala 37:23]
  wire [4:0] hazardu_io_rs2IDEX; // @[riscv.scala 37:23]
  wire  hazardu_io_regEnMEMWB; // @[riscv.scala 37:23]
  wire [4:0] hazardu_io_rdMEMWB; // @[riscv.scala 37:23]
  wire  hazardu_io_regEnWBEND; // @[riscv.scala 37:23]
  wire [4:0] hazardu_io_rdWBEND; // @[riscv.scala 37:23]
  wire [1:0] hazardu_io_forwardA; // @[riscv.scala 37:23]
  wire [1:0] hazardu_io_forwardB; // @[riscv.scala 37:23]
  wire [1:0] hazardu_io_forwardC; // @[riscv.scala 37:23]
  wire [4:0] hazardu_io_rs1IFID; // @[riscv.scala 37:23]
  wire [4:0] hazardu_io_rs2IFID; // @[riscv.scala 37:23]
  wire [4:0] hazardu_io_rdIDEX; // @[riscv.scala 37:23]
  wire [1:0] hazardu_io_resSrc; // @[riscv.scala 37:23]
  wire  hazardu_io_loadHazard; // @[riscv.scala 37:23]
  wire  preBranchIns_clock; // @[riscv.scala 38:28]
  wire  preBranchIns_reset; // @[riscv.scala 38:28]
  wire  preBranchIns_io_exjump; // @[riscv.scala 38:28]
  wire [31:0] preBranchIns_io_ifpc; // @[riscv.scala 38:28]
  wire [31:0] preBranchIns_io_expc; // @[riscv.scala 38:28]
  wire [31:0] preBranchIns_io_exdpc; // @[riscv.scala 38:28]
  wire [31:0] preBranchIns_io_ifdnpc; // @[riscv.scala 38:28]
  wire  preBranchIns_io_ifjump; // @[riscv.scala 38:28]
  wire  preBranchIns_block23_0; // @[riscv.scala 38:28]
  wire  preBranchIns_block1_0; // @[riscv.scala 38:28]
  wire [31:0] memVGenInst_io_inst; // @[riscv.scala 62:28]
  wire  memVGenInst_io_valid; // @[riscv.scala 62:28]
  wire [31:0] ctrl_io_inst; // @[riscv.scala 67:20]
  wire [1:0] ctrl_io_CtrlS_AluSrc1; // @[riscv.scala 67:20]
  wire [1:0] ctrl_io_CtrlS_AluSrc2; // @[riscv.scala 67:20]
  wire [4:0] ctrl_io_CtrlS_ALUCtrl; // @[riscv.scala 67:20]
  wire  ctrl_io_CtrlS_memWriteM; // @[riscv.scala 67:20]
  wire [7:0] ctrl_io_CtrlS_memWriteMask; // @[riscv.scala 67:20]
  wire [2:0] ctrl_io_CtrlS_memReadNum; // @[riscv.scala 67:20]
  wire  ctrl_io_CtrlS_dnpcSrc; // @[riscv.scala 67:20]
  wire  ctrl_io_CtrlS_jump; // @[riscv.scala 67:20]
  wire  ctrl_io_CtrlS_branch; // @[riscv.scala 67:20]
  wire  ctrl_io_CtrlS_regEn; // @[riscv.scala 67:20]
  wire [1:0] ctrl_io_CtrlS_ResultSrc; // @[riscv.scala 67:20]
  wire  ctrl_io_CtrlS_fencei; // @[riscv.scala 67:20]
  wire [31:0] csrCtrl_io_inst; // @[riscv.scala 68:23]
  wire  csrCtrl_io_CSRCtrlIf_csrrwen; // @[riscv.scala 68:23]
  wire  csrCtrl_io_CSRCtrlIf_csrswen; // @[riscv.scala 68:23]
  wire  csrCtrl_io_CSRCtrlIf_csrrsien; // @[riscv.scala 68:23]
  wire  csrCtrl_io_CSRCtrlIf_csrrcien; // @[riscv.scala 68:23]
  wire  csrCtrl_io_CSRCtrlIf_csrrcen; // @[riscv.scala 68:23]
  wire  csrCtrl_io_CSRCtrlIf_csrrwien; // @[riscv.scala 68:23]
  wire  csrCtrl_io_CSRCtrlIf_ecall; // @[riscv.scala 68:23]
  wire  csrCtrl_io_CSRCtrlIf_rfen; // @[riscv.scala 68:23]
  wire  csrCtrl_io_CSRCtrlIf_mepc2pc; // @[riscv.scala 68:23]
  wire  difftest_v; // @[riscv.scala 402:26]
  wire  intrins_intr; // @[riscv.scala 404:25]
  wire  Ebpro_block; // @[riscv.scala 406:23]
  wire [31:0] Ebpro_inst; // @[riscv.scala 406:23]
  wire  skipinst_v; // @[riscv.scala 410:26]
  wire  block1_0 = exu_block1;
  wire  _T = ~block1_0; // @[riscv.scala 55:32]
  wire  _T_2 = ~blockDMA_0; // @[riscv.scala 55:43]
  wire  _T_4 = ~io_instIO_ready; // @[riscv.scala 59:23]
  wire  _T_5 = _T_4; // @[riscv.scala 59:20]
  wire  block2 = _T_4; // @[riscv.scala 58:20 riscv.scala 59:10]
  reg [281:0] pipEX2MEMReg; // @[Reg.scala 27:20]
  wire  pipEX2MEMWire_valid = pipEX2MEMReg[80]; // @[riscv.scala 264:44]
  wire  _T_182 = ~io_dataIO_ready; // @[riscv.scala 279:36]
  wire  _T_183 = pipEX2MEMWire_valid & _T_182; // @[riscv.scala 279:33]
  wire  block3 = _T_183; // @[riscv.scala 278:20 riscv.scala 279:10]
  wire  _T_184 = _T_5 | block3; // @[riscv.scala 284:21]
  wire  block23 = _T_184; // @[riscv.scala 283:23 riscv.scala 284:11]
  wire  _T_252 = block1_0 | block23; // @[riscv.scala 393:22]
  wire  pipBlock = _T_252 | blockDMA_0; // @[riscv.scala 393:32]
  wire  _T_10 = ~pipBlock; // @[riscv.scala 88:30]
  reg [431:0] _T_68; // @[Reg.scala 27:20]
  wire  pipID2ExWire_branch = _T_68[49]; // @[riscv.scala 166:41]
  wire  _T_227 = pipID2ExWire_branch & exu_io_brTake; // @[riscv.scala 347:49]
  wire  pipID2ExWire_jump = _T_68[50]; // @[riscv.scala 166:41]
  wire  _T_228 = _T_227 | pipID2ExWire_jump; // @[riscv.scala 347:67]
  reg [8:0] _T_110; // @[Reg.scala 27:20]
  wire  pipCSRRegWire_mepc2pc = _T_110[0]; // @[riscv.scala 218:41]
  wire  _T_229 = _T_228 | pipCSRRegWire_mepc2pc; // @[riscv.scala 347:88]
  wire  pipCSRRegWire_ecall = _T_110[2]; // @[riscv.scala 218:41]
  wire  dnpcTakenWithoutPreB = _T_229 | pipCSRRegWire_ecall; // @[riscv.scala 347:113]
  wire  _T_231 = ~dnpcTakenWithoutPreB; // @[riscv.scala 348:15]
  wire  pipID2ExWire_ifjump = _T_68[34]; // @[riscv.scala 166:41]
  wire  jump1 = _T_231 & pipID2ExWire_ifjump; // @[riscv.scala 348:37]
  wire [31:0] pipID2ExWire_ifdnpc = _T_68[33:2]; // @[riscv.scala 166:41]
  wire  _T_232 = exu_io_dnpc != pipID2ExWire_ifdnpc; // @[riscv.scala 349:52]
  wire  _T_233 = ~pipID2ExWire_ifjump; // @[riscv.scala 349:79]
  wire  _T_234 = _T_232 | _T_233; // @[riscv.scala 349:76]
  wire  jump2 = dnpcTakenWithoutPreB & _T_234; // @[riscv.scala 349:36]
  wire  _T_235 = jump1 | jump2; // @[riscv.scala 350:25]
  wire [31:0] pipID2ExWire_pc = _T_68[142:111]; // @[riscv.scala 166:41]
  wire  _T_236 = pipID2ExWire_pc != 32'h0; // @[riscv.scala 350:69]
  wire  _T_237 = intrTimeCnt_0 & _T_236; // @[riscv.scala 350:50]
  wire  _T_238 = _T_235 | _T_237; // @[riscv.scala 350:34]
  wire  pipID2ExWire_fencei = _T_68[35]; // @[riscv.scala 166:41]
  wire  pipFlashWire = _T_238 | pipID2ExWire_fencei; // @[riscv.scala 350:78]
  wire  _T_11 = pipFlashWire & _T_10; // @[riscv.scala 88:27]
  wire  _T_13 = _T_11 | reset; // @[riscv.scala 88:40]
  wire  _T_14 = ifu_io_pc != 32'h0; // @[riscv.scala 90:16]
  wire [129:0] _T_19 = {_T_14,ifu_io_instOut,ifu_io_pc,ifu_io_snpc,preBranchIns_io_ifjump,preBranchIns_io_ifdnpc}; // @[Cat.scala 29:58]
  wire  _T_20 = pipBlock | hazardu_io_loadHazard; // @[riscv.scala 96:24]
  wire  _T_21 = ~_T_20; // @[riscv.scala 96:13]
  reg [129:0] _T_22; // @[Reg.scala 27:20]
  wire [31:0] pipIF2IDWire_ifdnpc = _T_22[31:0]; // @[riscv.scala 98:41]
  wire  pipIF2IDWire_ifjump = _T_22[32]; // @[riscv.scala 98:41]
  wire [31:0] pipIF2IDWire_snpc = _T_22[64:33]; // @[riscv.scala 98:41]
  wire [31:0] pipIF2IDWire_pc = _T_22[96:65]; // @[riscv.scala 98:41]
  wire [31:0] pipIF2IDWire_inst = _T_22[128:97]; // @[riscv.scala 98:41]
  wire  pipIF2IDWire_cmd = _T_22[129]; // @[riscv.scala 98:41]
  wire  _T_31 = pipFlashWire | hazardu_io_loadHazard; // @[riscv.scala 133:28]
  wire  _T_33 = _T_31 & _T_10; // @[riscv.scala 133:54]
  wire  _T_35 = _T_33 | reset; // @[riscv.scala 133:67]
  wire [31:0] _T_36 = pipIF2IDWire_inst & 32'hfe00707f; // @[riscv.scala 161:25]
  wire  _T_37 = 32'hc00607b == _T_36; // @[riscv.scala 161:25]
  wire  _T_39 = 32'he00707b == _T_36; // @[riscv.scala 162:25]
  wire [45:0] _T_45 = {idu_io_rs1,idu_io_rs2,ctrl_io_CtrlS_fencei,pipIF2IDWire_ifjump,pipIF2IDWire_ifdnpc,_T_37,_T_39}; // @[Cat.scala 29:58]
  wire [60:0] _T_52 = {ctrl_io_CtrlS_memWriteMask,ctrl_io_CtrlS_memWriteM,ctrl_io_CtrlS_dnpcSrc,ctrl_io_CtrlS_jump,ctrl_io_CtrlS_branch,ctrl_io_CtrlS_regEn,ctrl_io_CtrlS_ResultSrc,_T_45}; // @[Cat.scala 29:58]
  wire [49:0] _T_58 = {pipIF2IDWire_snpc,idu_io_rdOut,ctrl_io_CtrlS_ALUCtrl,ctrl_io_CtrlS_AluSrc1,ctrl_io_CtrlS_AluSrc2,ctrl_io_CtrlS_memReadNum,memVGenInst_io_valid}; // @[Cat.scala 29:58]
  wire [431:0] _T_66 = {pipIF2IDWire_cmd,pipIF2IDWire_inst,idu_io_dataEx_imme,idu_io_dataEx_dOut1,idu_io_dataEx_dOut2,idu_io_dataEx_rdDout,pipIF2IDWire_pc,_T_58,_T_52}; // @[Cat.scala 29:58]
  wire  pipID2ExWire_dmaWR = _T_68[0]; // @[riscv.scala 166:41]
  wire  pipID2ExWire_dma = _T_68[1]; // @[riscv.scala 166:41]
  wire [1:0] pipID2ExWire_resultSrc = _T_68[47:46]; // @[riscv.scala 166:41]
  wire  pipID2ExWire_regEn = _T_68[48]; // @[riscv.scala 166:41]
  wire  pipID2ExWire_memWriteM = _T_68[52]; // @[riscv.scala 166:41]
  wire [7:0] pipID2ExWire_mask = _T_68[60:53]; // @[riscv.scala 166:41]
  wire  pipID2ExWire_valid = _T_68[61]; // @[riscv.scala 166:41]
  wire [2:0] pipID2ExWire_memReadNum = _T_68[64:62]; // @[riscv.scala 166:41]
  wire [4:0] pipID2ExWire_rd = _T_68[78:74]; // @[riscv.scala 166:41]
  wire [31:0] pipID2ExWire_snpc = _T_68[110:79]; // @[riscv.scala 166:41]
  wire [31:0] pipID2ExWire_inst = _T_68[430:399]; // @[riscv.scala 166:41]
  wire  pipID2ExWire_cmd = _T_68[431]; // @[riscv.scala 166:41]
  wire [8:0] _T_108 = {csrCtrl_io_CSRCtrlIf_csrrwen,csrCtrl_io_CSRCtrlIf_csrswen,csrCtrl_io_CSRCtrlIf_csrrsien,csrCtrl_io_CSRCtrlIf_csrrcien,csrCtrl_io_CSRCtrlIf_csrrcen,csrCtrl_io_CSRCtrlIf_csrrwien,csrCtrl_io_CSRCtrlIf_ecall,csrCtrl_io_CSRCtrlIf_rfen,csrCtrl_io_CSRCtrlIf_mepc2pc}; // @[Cat.scala 29:58]
  wire  pipCSRRegWire_rfen = _T_110[1]; // @[riscv.scala 218:41]
  wire  _T_124 = pipID2ExWire_regEn | pipCSRRegWire_rfen; // @[riscv.scala 254:21]
  wire  _T_69_dma = pipID2ExWire_dma; // @[riscv.scala 166:41 riscv.scala 166:41]
  wire  _T_69_dmaWR = pipID2ExWire_dmaWR; // @[riscv.scala 166:41 riscv.scala 166:41]
  wire  _T_127 = pipID2ExWire_dma | pipID2ExWire_dmaWR; // @[riscv.scala 259:22]
  wire [71:0] _T_135 = {pipID2ExWire_memWriteM,_T_124,pipID2ExWire_resultSrc,pipID2ExWire_pc,pipID2ExWire_fencei,_T_237,_T_127,exu_io_dnpc,dnpcTakenWithoutPreB}; // @[Cat.scala 29:58]
  wire [281:0] _T_144 = {pipID2ExWire_cmd,pipID2ExWire_inst,exu_io_dataOut_ALUResOut,exu_io_dataOut_wdata,pipID2ExWire_snpc,pipID2ExWire_rd,pipID2ExWire_memReadNum,pipID2ExWire_valid,pipID2ExWire_mask,_T_135}; // @[Cat.scala 29:58]
  wire  pipEX2MEMWire_skip = pipEX2MEMReg[33]; // @[riscv.scala 264:44]
  wire  pipEX2MEMWire_intr = pipEX2MEMReg[34]; // @[riscv.scala 264:44]
  wire  pipEX2MEMWire_fencei = pipEX2MEMReg[35]; // @[riscv.scala 264:44]
  wire [31:0] pipEX2MEMWire_pc = pipEX2MEMReg[67:36]; // @[riscv.scala 264:44]
  wire [1:0] pipEX2MEMWire_ResultSrc = pipEX2MEMReg[69:68]; // @[riscv.scala 264:44]
  wire  pipEX2MEMWire_regEn = pipEX2MEMReg[70]; // @[riscv.scala 264:44]
  wire [7:0] pipEX2MEMWire_mask = pipEX2MEMReg[79:72]; // @[riscv.scala 264:44]
  wire [2:0] pipEX2MEMWire_memReadNum = pipEX2MEMReg[83:81]; // @[riscv.scala 264:44]
  wire [4:0] pipEX2MEMWire_rd = pipEX2MEMReg[88:84]; // @[riscv.scala 264:44]
  wire [31:0] pipEX2MEMWire_snpc = pipEX2MEMReg[120:89]; // @[riscv.scala 264:44]
  wire [63:0] pipEX2MEMWire_writeDataM = pipEX2MEMReg[184:121]; // @[riscv.scala 264:44]
  wire [63:0] pipEX2MEMWire_ALURes = pipEX2MEMReg[248:185]; // @[riscv.scala 264:44]
  wire [31:0] pipEX2MEMWire_inst = pipEX2MEMReg[280:249]; // @[riscv.scala 264:44]
  wire  pipEX2MEMWire_cmd = pipEX2MEMReg[281]; // @[riscv.scala 264:44]
  wire [14:0] _GEN_7 = {{7'd0}, pipEX2MEMWire_mask}; // @[riscv.scala 267:40]
  wire [14:0] _T_167 = _GEN_7 << pipEX2MEMWire_ALURes[2:0]; // @[riscv.scala 267:40]
  wire [3:0] _GEN_8 = {{1'd0}, pipEX2MEMWire_ALURes[2:0]}; // @[riscv.scala 272:78]
  wire [6:0] _T_170 = _GEN_8 * 4'h8; // @[riscv.scala 272:78]
  wire [190:0] _GEN_9 = {{127'd0}, pipEX2MEMWire_writeDataM}; // @[riscv.scala 272:50]
  wire [190:0] _T_171 = _GEN_9 << _T_170; // @[riscv.scala 272:50]
  wire  _T_173 = pipEX2MEMWire_valid & _T; // @[riscv.scala 273:42]
  wire  _T_176 = pipEX2MEMWire_ResultSrc == 2'h0; // @[riscv.scala 274:49]
  wire  _T_178 = pipEX2MEMWire_ALURes < 64'h80000000; // @[riscv.scala 276:59]
  wire  _T_179 = pipEX2MEMWire_ALURes > 64'h8fffffff; // @[riscv.scala 276:95]
  wire  _T_180 = _T_178 | _T_179; // @[riscv.scala 276:71]
  wire  _T_181 = pipEX2MEMWire_valid & _T_180; // @[riscv.scala 276:34]
  wire  skip = _T_181 | pipEX2MEMWire_fencei; // @[riscv.scala 276:109]
  wire  jud = pipEX2MEMWire_pc == 32'h0; // @[riscv.scala 289:29]
  wire  _T_185 = skip | pipEX2MEMWire_skip; // @[riscv.scala 302:10]
  reg [173:0] pipMEM2WBReg; // @[Reg.scala 27:20]
  wire [31:0] pipMEM2WBWire_pc = pipMEM2WBReg[33:2]; // @[riscv.scala 304:44]
  wire [31:0] _T_210 = pipMEM2WBWire_pc + 32'h4; // @[riscv.scala 305:42]
  wire [31:0] npcsend = jud ? _T_210 : pipEX2MEMWire_pc; // @[riscv.scala 305:17]
  wire [36:0] _T_189 = {pipEX2MEMWire_regEn,pipEX2MEMWire_ResultSrc,npcsend,pipEX2MEMWire_intr,_T_185}; // @[Cat.scala 29:58]
  wire [173:0] _T_195 = {pipEX2MEMWire_cmd,pipEX2MEMWire_inst,pipEX2MEMWire_ALURes,pipEX2MEMWire_rd,pipEX2MEMWire_snpc,pipEX2MEMWire_memReadNum,_T_189}; // @[Cat.scala 29:58]
  wire  pipMEM2WBWire_intr = pipMEM2WBReg[1]; // @[riscv.scala 304:44]
  wire  pipMEM2WBWire_regEn = pipMEM2WBReg[36]; // @[riscv.scala 304:44]
  wire [4:0] pipMEM2WBWire_rd = pipMEM2WBReg[76:72]; // @[riscv.scala 304:44]
  wire [63:0] pipMEM2WBWire_ALURes = pipMEM2WBReg[140:77]; // @[riscv.scala 304:44]
  wire [31:0] pipMEM2WBWire_inst = pipMEM2WBReg[172:141]; // @[riscv.scala 304:44]
  wire  pipMEM2WBWire_cmd = pipMEM2WBReg[173]; // @[riscv.scala 304:44]
  reg [63:0] _T_213; // @[Reg.scala 27:20]
  wire [3:0] _GEN_10 = {{1'd0}, pipMEM2WBWire_ALURes[2:0]}; // @[riscv.scala 313:100]
  wire [6:0] _T_215 = _GEN_10 * 4'h8; // @[riscv.scala 313:100]
  wire [69:0] _T_219 = {pipMEM2WBWire_rd,pipMEM2WBWire_regEn,pipMEM2WBWire_inst,pipMEM2WBWire_pc}; // @[Cat.scala 29:58]
  reg [69:0] _T_221; // @[Reg.scala 27:20]
  wire [31:0] _T_248 = jump2 ? exu_io_dnpc : preBranchIns_io_ifdnpc; // @[riscv.scala 362:12]
  wire [31:0] _T_249 = jump1 ? pipID2ExWire_snpc : _T_248; // @[riscv.scala 359:10]
  wire [31:0] _T_250 = pipID2ExWire_fencei ? pipID2ExWire_snpc : _T_249; // @[riscv.scala 356:8]
  wire  _T_254 = ~intrTimeCnt_0; // @[riscv.scala 396:36]
  wire  _T_255 = pipID2ExWire_fencei & _T_254; // @[riscv.scala 396:33]
  wire  _T_257 = _T_255 & _T_10; // @[riscv.scala 396:49]
  wire  hazardPCBlock = hazardu_io_loadHazard; // @[riscv.scala 389:27 riscv.scala 390:17]
  wire  _T_99 = pipID2ExWire_dma; // @[riscv.scala 168:21 riscv.scala 169:11]
  wire  _T_100 = pipID2ExWire_dmaWR; // @[riscv.scala 172:23 riscv.scala 173:13]
  wire  fencei = _T_257; // @[riscv.scala 395:20 riscv.scala 396:10]
  iFetch ifu ( // @[riscv.scala 34:19]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_instIn(ifu_io_instIn),
    .io_instOut(ifu_io_instOut),
    .io_pc(ifu_io_pc),
    .io_snpc(ifu_io_snpc),
    .io_dnpc(ifu_io_dnpc),
    .io_jump(ifu_io_jump),
    .intrTimeCnt_0(ifu_intrTimeCnt_0),
    .hazardPCBlock_0(ifu_hazardPCBlock_0),
    .blockDMA_0(ifu_blockDMA_0),
    .block23_0(ifu_block23_0),
    .block1_0(ifu_block1_0)
  );
  iDecode idu ( // @[riscv.scala 35:19]
    .clock(idu_clock),
    .reset(idu_reset),
    .io_pc(idu_io_pc),
    .io_inst(idu_io_inst),
    .io_regEn(idu_io_regEn),
    .io_dataEx_imme(idu_io_dataEx_imme),
    .io_dataEx_dOut1(idu_io_dataEx_dOut1),
    .io_dataEx_dOut2(idu_io_dataEx_dOut2),
    .io_dataEx_dIn(idu_io_dataEx_dIn),
    .io_dataEx_rdDout(idu_io_dataEx_rdDout),
    .io_rdOut(idu_io_rdOut),
    .io_rdIn(idu_io_rdIn),
    .io_rs1(idu_io_rs1),
    .io_rs2(idu_io_rs2),
    .io_dOutWB(idu_io_dOutWB),
    .blockDMA(idu_blockDMA),
    .block23(idu_block23),
    .block1(idu_block1)
  );
  execute exu ( // @[riscv.scala 36:19]
    .clock(exu_clock),
    .reset(exu_reset),
    .io_AluSrc1(exu_io_AluSrc1),
    .io_AluSrc2(exu_io_AluSrc2),
    .io_ALUCtrl(exu_io_ALUCtrl),
    .io_dnpcSrc(exu_io_dnpcSrc),
    .io_ResultSrc(exu_io_ResultSrc),
    .io_memReadNum(exu_io_memReadNum),
    .io_dataId_imme(exu_io_dataId_imme),
    .io_dataId_dOut1(exu_io_dataId_dOut1),
    .io_dataId_dOut2(exu_io_dataId_dOut2),
    .io_dataId_dIn(exu_io_dataId_dIn),
    .io_dataId_rdDout(exu_io_dataId_rdDout),
    .io_dataOut_ALUResOut(exu_io_dataOut_ALUResOut),
    .io_dataOut_wdata(exu_io_dataOut_wdata),
    .io_dataOut_rdata(exu_io_dataOut_rdata),
    .io_brTake(exu_io_brTake),
    .io_pc(exu_io_pc),
    .io_snpc(exu_io_snpc),
    .io_dnpc(exu_io_dnpc),
    .io_CSRCtrlIf_csrrwen(exu_io_CSRCtrlIf_csrrwen),
    .io_CSRCtrlIf_csrswen(exu_io_CSRCtrlIf_csrswen),
    .io_CSRCtrlIf_csrrsien(exu_io_CSRCtrlIf_csrrsien),
    .io_CSRCtrlIf_csrrcien(exu_io_CSRCtrlIf_csrrcien),
    .io_CSRCtrlIf_csrrcen(exu_io_CSRCtrlIf_csrrcen),
    .io_CSRCtrlIf_csrrwien(exu_io_CSRCtrlIf_csrrwien),
    .io_CSRCtrlIf_ecall(exu_io_CSRCtrlIf_ecall),
    .io_CSRCtrlIf_rfen(exu_io_CSRCtrlIf_rfen),
    .io_CSRCtrlIf_mepc2pc(exu_io_CSRCtrlIf_mepc2pc),
    .io_uimm(exu_io_uimm),
    .io_aluResIn(exu_io_aluResIn),
    .io_forwardA(exu_io_forwardA),
    .io_forwardB(exu_io_forwardB),
    .io_forwardC(exu_io_forwardC),
    .io_aluRes1(exu_io_aluRes1),
    .io_aluRes3(exu_io_aluRes3),
    .intrTimeCnt_0(exu_intrTimeCnt_0),
    .startTimeCnt(exu_startTimeCnt),
    .dmaCtrl_0(exu_dmaCtrl_0),
    .blockDMA(exu_blockDMA),
    .block23(exu_block23),
    .block1(exu_block1)
  );
  hazard hazardu ( // @[riscv.scala 37:23]
    .io_regEnEXMEM(hazardu_io_regEnEXMEM),
    .io_rdEXMEM(hazardu_io_rdEXMEM),
    .io_rs1IDEX(hazardu_io_rs1IDEX),
    .io_rs2IDEX(hazardu_io_rs2IDEX),
    .io_regEnMEMWB(hazardu_io_regEnMEMWB),
    .io_rdMEMWB(hazardu_io_rdMEMWB),
    .io_regEnWBEND(hazardu_io_regEnWBEND),
    .io_rdWBEND(hazardu_io_rdWBEND),
    .io_forwardA(hazardu_io_forwardA),
    .io_forwardB(hazardu_io_forwardB),
    .io_forwardC(hazardu_io_forwardC),
    .io_rs1IFID(hazardu_io_rs1IFID),
    .io_rs2IFID(hazardu_io_rs2IFID),
    .io_rdIDEX(hazardu_io_rdIDEX),
    .io_resSrc(hazardu_io_resSrc),
    .io_loadHazard(hazardu_io_loadHazard)
  );
  preBranch preBranchIns ( // @[riscv.scala 38:28]
    .clock(preBranchIns_clock),
    .reset(preBranchIns_reset),
    .io_exjump(preBranchIns_io_exjump),
    .io_ifpc(preBranchIns_io_ifpc),
    .io_expc(preBranchIns_io_expc),
    .io_exdpc(preBranchIns_io_exdpc),
    .io_ifdnpc(preBranchIns_io_ifdnpc),
    .io_ifjump(preBranchIns_io_ifjump),
    .block23_0(preBranchIns_block23_0),
    .block1_0(preBranchIns_block1_0)
  );
  memVGen memVGenInst ( // @[riscv.scala 62:28]
    .io_inst(memVGenInst_io_inst),
    .io_valid(memVGenInst_io_valid)
  );
  CtrlUnit ctrl ( // @[riscv.scala 67:20]
    .io_inst(ctrl_io_inst),
    .io_CtrlS_AluSrc1(ctrl_io_CtrlS_AluSrc1),
    .io_CtrlS_AluSrc2(ctrl_io_CtrlS_AluSrc2),
    .io_CtrlS_ALUCtrl(ctrl_io_CtrlS_ALUCtrl),
    .io_CtrlS_memWriteM(ctrl_io_CtrlS_memWriteM),
    .io_CtrlS_memWriteMask(ctrl_io_CtrlS_memWriteMask),
    .io_CtrlS_memReadNum(ctrl_io_CtrlS_memReadNum),
    .io_CtrlS_dnpcSrc(ctrl_io_CtrlS_dnpcSrc),
    .io_CtrlS_jump(ctrl_io_CtrlS_jump),
    .io_CtrlS_branch(ctrl_io_CtrlS_branch),
    .io_CtrlS_regEn(ctrl_io_CtrlS_regEn),
    .io_CtrlS_ResultSrc(ctrl_io_CtrlS_ResultSrc),
    .io_CtrlS_fencei(ctrl_io_CtrlS_fencei)
  );
  csrCtrl csrCtrl ( // @[riscv.scala 68:23]
    .io_inst(csrCtrl_io_inst),
    .io_CSRCtrlIf_csrrwen(csrCtrl_io_CSRCtrlIf_csrrwen),
    .io_CSRCtrlIf_csrswen(csrCtrl_io_CSRCtrlIf_csrswen),
    .io_CSRCtrlIf_csrrsien(csrCtrl_io_CSRCtrlIf_csrrsien),
    .io_CSRCtrlIf_csrrcien(csrCtrl_io_CSRCtrlIf_csrrcien),
    .io_CSRCtrlIf_csrrcen(csrCtrl_io_CSRCtrlIf_csrrcen),
    .io_CSRCtrlIf_csrrwien(csrCtrl_io_CSRCtrlIf_csrrwien),
    .io_CSRCtrlIf_ecall(csrCtrl_io_CSRCtrlIf_ecall),
    .io_CSRCtrlIf_rfen(csrCtrl_io_CSRCtrlIf_rfen),
    .io_CSRCtrlIf_mepc2pc(csrCtrl_io_CSRCtrlIf_mepc2pc)
  );
  difftest difftest ( // @[riscv.scala 402:26]
    .v(difftest_v)
  );
  intr intrins ( // @[riscv.scala 404:25]
    .intr(intrins_intr)
  );
  ebProbe Ebpro ( // @[riscv.scala 406:23]
    .block(Ebpro_block),
    .inst(Ebpro_inst)
  );
  skip skipinst ( // @[riscv.scala 410:26]
    .v(skipinst_v)
  );
  assign io_instIO_valid = _T & _T_2; // @[riscv.scala 55:19]
  assign io_instIO_addr = ifu_io_pc; // @[riscv.scala 81:18]
  assign io_dataIO_valid = _T_173 & _T_2; // @[riscv.scala 273:19]
  assign io_dataIO_data_write = _T_171[63:0]; // @[riscv.scala 272:23]
  assign io_dataIO_wen = pipEX2MEMReg[71]; // @[riscv.scala 268:17]
  assign io_dataIO_addr = pipEX2MEMWire_ALURes[31:0]; // @[riscv.scala 270:18]
  assign io_dataIO_rsize = pipEX2MEMWire_memReadNum[1:0]; // @[riscv.scala 271:19]
  assign io_dataIO_mask = _T_167[7:0]; // @[riscv.scala 267:18]
  assign _T_99_0 = _T_69_dma;
  assign _T_100_0 = _T_69_dmaWR;
  assign startTimeCnt = exu_startTimeCnt;
  assign block3_0 = block3;
  assign dmaCtrl = exu_dmaCtrl_0;
  assign block2_0 = _T_5;
  assign fencei_0 = fencei;
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_instIn = ifu_io_pc[2] ? io_instIO_data_read[63:32] : io_instIO_data_read[31:0]; // @[riscv.scala 80:17]
  assign ifu_io_dnpc = _T_237 ? exu_io_dnpc : _T_250; // @[riscv.scala 353:15]
  assign ifu_io_jump = pipFlashWire | preBranchIns_io_ifjump; // @[riscv.scala 352:15]
  assign ifu_intrTimeCnt_0 = intrTimeCnt_0;
  assign ifu_hazardPCBlock_0 = hazardPCBlock;
  assign ifu_blockDMA_0 = blockDMA_0;
  assign ifu_block23_0 = block23;
  assign ifu_block1_0 = exu_block1;
  assign idu_clock = clock;
  assign idu_reset = reset;
  assign idu_io_pc = pipMEM2WBReg[33:2]; // @[riscv.scala 316:13]
  assign idu_io_inst = _T_22[128:97]; // @[riscv.scala 103:17]
  assign idu_io_regEn = pipMEM2WBReg[36]; // @[riscv.scala 310:16]
  assign idu_io_dataEx_dIn = exu_io_dataId_dIn; // @[riscv.scala 314:21]
  assign idu_io_rdIn = pipMEM2WBReg[76:72]; // @[riscv.scala 307:15]
  assign idu_blockDMA = blockDMA_0;
  assign idu_block23 = block23;
  assign idu_block1 = exu_block1;
  assign exu_clock = clock;
  assign exu_reset = reset;
  assign exu_io_AluSrc1 = _T_68[68:67]; // @[riscv.scala 185:20]
  assign exu_io_AluSrc2 = _T_68[66:65]; // @[riscv.scala 186:20]
  assign exu_io_ALUCtrl = _T_68[73:69]; // @[riscv.scala 184:19]
  assign exu_io_dnpcSrc = _T_68[51]; // @[riscv.scala 191:20]
  assign exu_io_ResultSrc = pipMEM2WBReg[35:34]; // @[riscv.scala 311:20]
  assign exu_io_memReadNum = pipMEM2WBReg[39:37]; // @[riscv.scala 309:21]
  assign exu_io_dataId_imme = _T_68[398:335]; // @[riscv.scala 177:24]
  assign exu_io_dataId_dOut1 = _T_68[334:271]; // @[riscv.scala 178:25]
  assign exu_io_dataId_dOut2 = _T_68[270:207]; // @[riscv.scala 179:25]
  assign exu_io_dataId_rdDout = _T_68[206:143]; // @[riscv.scala 180:26]
  assign exu_io_dataOut_rdata = _T_213 >> _T_215; // @[riscv.scala 313:24]
  assign exu_io_pc = _T_68[142:111]; // @[riscv.scala 181:15]
  assign exu_io_snpc = pipMEM2WBReg[71:40]; // @[riscv.scala 308:15]
  assign exu_io_CSRCtrlIf_csrrwen = _T_110[8]; // @[riscv.scala 219:30]
  assign exu_io_CSRCtrlIf_csrswen = _T_110[7]; // @[riscv.scala 220:30]
  assign exu_io_CSRCtrlIf_csrrsien = _T_110[6]; // @[riscv.scala 221:31]
  assign exu_io_CSRCtrlIf_csrrcien = _T_110[5]; // @[riscv.scala 222:31]
  assign exu_io_CSRCtrlIf_csrrcen = _T_110[4]; // @[riscv.scala 223:30]
  assign exu_io_CSRCtrlIf_csrrwien = _T_110[3]; // @[riscv.scala 224:31]
  assign exu_io_CSRCtrlIf_ecall = _T_110[2]; // @[riscv.scala 225:28]
  assign exu_io_CSRCtrlIf_rfen = _T_110[1]; // @[riscv.scala 226:27]
  assign exu_io_CSRCtrlIf_mepc2pc = _T_110[0]; // @[riscv.scala 228:30]
  assign exu_io_uimm = _T_68[45:41]; // @[riscv.scala 229:17]
  assign exu_io_aluResIn = pipMEM2WBReg[140:77]; // @[riscv.scala 306:19]
  assign exu_io_forwardA = hazardu_io_forwardA; // @[riscv.scala 379:19]
  assign exu_io_forwardB = hazardu_io_forwardB; // @[riscv.scala 380:19]
  assign exu_io_forwardC = hazardu_io_forwardC; // @[riscv.scala 381:19]
  assign exu_io_aluRes1 = _T_176 ? pipEX2MEMWire_ALURes : {{32'd0}, pipEX2MEMWire_snpc}; // @[riscv.scala 274:18]
  assign exu_io_aluRes3 = idu_io_dOutWB; // @[riscv.scala 343:18]
  assign exu_intrTimeCnt_0 = intrTimeCnt_0;
  assign exu_blockDMA = blockDMA_0;
  assign exu_block23 = block23;
  assign hazardu_io_regEnEXMEM = pipEX2MEMReg[70]; // @[riscv.scala 372:25]
  assign hazardu_io_rdEXMEM = pipEX2MEMReg[88:84]; // @[riscv.scala 373:22]
  assign hazardu_io_rs1IDEX = _T_68[45:41]; // @[riscv.scala 198:24]
  assign hazardu_io_rs2IDEX = _T_68[40:36]; // @[riscv.scala 199:24]
  assign hazardu_io_regEnMEMWB = pipMEM2WBReg[36]; // @[riscv.scala 374:25]
  assign hazardu_io_rdMEMWB = pipMEM2WBReg[76:72]; // @[riscv.scala 375:22]
  assign hazardu_io_regEnWBEND = _T_221[64]; // @[riscv.scala 376:25]
  assign hazardu_io_rdWBEND = _T_221[69:65]; // @[riscv.scala 377:22]
  assign hazardu_io_rs1IFID = idu_io_rs1; // @[riscv.scala 384:22]
  assign hazardu_io_rs2IFID = idu_io_rs2; // @[riscv.scala 385:22]
  assign hazardu_io_rdIDEX = _T_68[78:74]; // @[riscv.scala 386:21]
  assign hazardu_io_resSrc = _T_68[47:46]; // @[riscv.scala 387:21]
  assign preBranchIns_clock = clock;
  assign preBranchIns_reset = reset;
  assign preBranchIns_io_exjump = pipEX2MEMReg[0]; // @[riscv.scala 417:28]
  assign preBranchIns_io_ifpc = ifu_io_pc; // @[riscv.scala 416:26]
  assign preBranchIns_io_expc = pipEX2MEMReg[67:36]; // @[riscv.scala 418:26]
  assign preBranchIns_io_exdpc = pipEX2MEMReg[32:1]; // @[riscv.scala 419:27]
  assign preBranchIns_block23_0 = block23;
  assign preBranchIns_block1_0 = exu_block1;
  assign memVGenInst_io_inst = _T_22[128:97]; // @[riscv.scala 100:25]
  assign ctrl_io_inst = _T_22[128:97]; // @[riscv.scala 102:18]
  assign csrCtrl_io_inst = _T_22[128:97]; // @[riscv.scala 101:21]
  assign difftest_v = pipMEM2WBWire_cmd & _T_10; // @[riscv.scala 403:19]
  assign intrins_intr = pipMEM2WBWire_intr & _T_10; // @[riscv.scala 405:21]
  assign Ebpro_block = _T_252 | blockDMA_0; // @[riscv.scala 408:20]
  assign Ebpro_inst = pipMEM2WBReg[172:141]; // @[riscv.scala 407:19]
  assign skipinst_v = pipMEM2WBReg[0]; // @[riscv.scala 411:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {9{`RANDOM}};
  pipEX2MEMReg = _RAND_0[281:0];
  _RAND_1 = {14{`RANDOM}};
  _T_68 = _RAND_1[431:0];
  _RAND_2 = {1{`RANDOM}};
  _T_110 = _RAND_2[8:0];
  _RAND_3 = {5{`RANDOM}};
  _T_22 = _RAND_3[129:0];
  _RAND_4 = {6{`RANDOM}};
  pipMEM2WBReg = _RAND_4[173:0];
  _RAND_5 = {2{`RANDOM}};
  _T_213 = _RAND_5[63:0];
  _RAND_6 = {3{`RANDOM}};
  _T_221 = _RAND_6[69:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pipEX2MEMReg <= 282'h0;
    end else if (_T_10) begin
      if (_T_237) begin
        pipEX2MEMReg <= 282'h1;
      end else begin
        pipEX2MEMReg <= _T_144;
      end
    end
    if (_T_35) begin
      _T_68 <= 432'h0;
    end else if (_T_10) begin
      _T_68 <= _T_66;
    end
    if (_T_35) begin
      _T_110 <= 9'h0;
    end else if (_T_10) begin
      _T_110 <= _T_108;
    end
    if (_T_13) begin
      _T_22 <= 130'h0;
    end else if (_T_21) begin
      _T_22 <= _T_19;
    end
    if (reset) begin
      pipMEM2WBReg <= 174'h0;
    end else if (_T_10) begin
      pipMEM2WBReg <= _T_195;
    end
    if (reset) begin
      _T_213 <= 64'h0;
    end else if (_T_10) begin
      _T_213 <= io_dataIO_data_read;
    end
    if (reset) begin
      _T_221 <= 70'h0;
    end else if (_T_10) begin
      _T_221 <= _T_219;
    end
  end
endmodule
module Icache(
  input          clock,
  input          reset,
  output         io_cacheOut_ar_valid_o,
  output [31:0]  io_cacheOut_ar_addr_o,
  output [7:0]   io_cacheOut_ar_len_o,
  input          io_cacheOut_r_valid_i,
  input  [63:0]  io_cacheOut_r_data_i,
  input          io_cacheOut_r_last_i,
  output [31:0]  io_cacheOut_w_addr_o,
  input          io_cacheIn_valid,
  output         io_cacheIn_ready,
  output [63:0]  io_cacheIn_data_read,
  input  [31:0]  io_cacheIn_addr,
  output         io_SRAMIO_0_cen,
  output         io_SRAMIO_0_wen,
  output [127:0] io_SRAMIO_0_wdata,
  output [5:0]   io_SRAMIO_0_addr,
  output [127:0] io_SRAMIO_0_wmask,
  input  [127:0] io_SRAMIO_0_rdata,
  output         io_SRAMIO_1_cen,
  output         io_SRAMIO_1_wen,
  output [127:0] io_SRAMIO_1_wdata,
  output [5:0]   io_SRAMIO_1_addr,
  output [127:0] io_SRAMIO_1_wmask,
  input  [127:0] io_SRAMIO_1_rdata,
  output         io_SRAMIO_2_cen,
  output         io_SRAMIO_2_wen,
  output [127:0] io_SRAMIO_2_wdata,
  output [5:0]   io_SRAMIO_2_addr,
  output [127:0] io_SRAMIO_2_wmask,
  input  [127:0] io_SRAMIO_2_rdata,
  output         io_SRAMIO_3_cen,
  output         io_SRAMIO_3_wen,
  output [127:0] io_SRAMIO_3_wdata,
  output [5:0]   io_SRAMIO_3_addr,
  output [127:0] io_SRAMIO_3_wmask,
  input  [127:0] io_SRAMIO_3_rdata,
  input          io_block,
  input          updataICache
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] _T_4; // @[Cache.scala 389:27]
  wire  _T_273 = 6'h3f == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_4289; // @[Reg.scala 27:20]
  wire  _T_271 = 6'h3e == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_4228; // @[Reg.scala 27:20]
  wire  _T_269 = 6'h3d == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_4167; // @[Reg.scala 27:20]
  wire  _T_267 = 6'h3c == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_4106; // @[Reg.scala 27:20]
  wire  _T_265 = 6'h3b == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_4045; // @[Reg.scala 27:20]
  wire  _T_263 = 6'h3a == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3984; // @[Reg.scala 27:20]
  wire  _T_261 = 6'h39 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3923; // @[Reg.scala 27:20]
  wire  _T_259 = 6'h38 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3862; // @[Reg.scala 27:20]
  wire  _T_257 = 6'h37 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3801; // @[Reg.scala 27:20]
  wire  _T_255 = 6'h36 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3740; // @[Reg.scala 27:20]
  wire  _T_253 = 6'h35 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3679; // @[Reg.scala 27:20]
  wire  _T_251 = 6'h34 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3618; // @[Reg.scala 27:20]
  wire  _T_249 = 6'h33 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3557; // @[Reg.scala 27:20]
  wire  _T_247 = 6'h32 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3496; // @[Reg.scala 27:20]
  wire  _T_245 = 6'h31 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3435; // @[Reg.scala 27:20]
  wire  _T_243 = 6'h30 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3374; // @[Reg.scala 27:20]
  wire  _T_241 = 6'h2f == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3313; // @[Reg.scala 27:20]
  wire  _T_239 = 6'h2e == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3252; // @[Reg.scala 27:20]
  wire  _T_237 = 6'h2d == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3191; // @[Reg.scala 27:20]
  wire  _T_235 = 6'h2c == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3130; // @[Reg.scala 27:20]
  wire  _T_233 = 6'h2b == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3069; // @[Reg.scala 27:20]
  wire  _T_231 = 6'h2a == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3008; // @[Reg.scala 27:20]
  wire  _T_229 = 6'h29 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2947; // @[Reg.scala 27:20]
  wire  _T_227 = 6'h28 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2886; // @[Reg.scala 27:20]
  wire  _T_225 = 6'h27 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2825; // @[Reg.scala 27:20]
  wire  _T_223 = 6'h26 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2764; // @[Reg.scala 27:20]
  wire  _T_221 = 6'h25 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2703; // @[Reg.scala 27:20]
  wire  _T_219 = 6'h24 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2642; // @[Reg.scala 27:20]
  wire  _T_217 = 6'h23 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2581; // @[Reg.scala 27:20]
  wire  _T_215 = 6'h22 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2520; // @[Reg.scala 27:20]
  wire  _T_213 = 6'h21 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2459; // @[Reg.scala 27:20]
  wire  _T_211 = 6'h20 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2398; // @[Reg.scala 27:20]
  wire  _T_209 = 6'h1f == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2337; // @[Reg.scala 27:20]
  wire  _T_207 = 6'h1e == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2276; // @[Reg.scala 27:20]
  wire  _T_205 = 6'h1d == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2215; // @[Reg.scala 27:20]
  wire  _T_203 = 6'h1c == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2154; // @[Reg.scala 27:20]
  wire  _T_201 = 6'h1b == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2093; // @[Reg.scala 27:20]
  wire  _T_199 = 6'h1a == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2032; // @[Reg.scala 27:20]
  wire  _T_197 = 6'h19 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1971; // @[Reg.scala 27:20]
  wire  _T_195 = 6'h18 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1910; // @[Reg.scala 27:20]
  wire  _T_193 = 6'h17 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1849; // @[Reg.scala 27:20]
  wire  _T_191 = 6'h16 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1788; // @[Reg.scala 27:20]
  wire  _T_189 = 6'h15 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1727; // @[Reg.scala 27:20]
  wire  _T_187 = 6'h14 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1666; // @[Reg.scala 27:20]
  wire  _T_185 = 6'h13 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1605; // @[Reg.scala 27:20]
  wire  _T_183 = 6'h12 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1544; // @[Reg.scala 27:20]
  wire  _T_181 = 6'h11 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1483; // @[Reg.scala 27:20]
  wire  _T_179 = 6'h10 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1422; // @[Reg.scala 27:20]
  wire  _T_177 = 6'hf == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1361; // @[Reg.scala 27:20]
  wire  _T_175 = 6'he == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1300; // @[Reg.scala 27:20]
  wire  _T_173 = 6'hd == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1239; // @[Reg.scala 27:20]
  wire  _T_171 = 6'hc == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1178; // @[Reg.scala 27:20]
  wire  _T_169 = 6'hb == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1117; // @[Reg.scala 27:20]
  wire  _T_167 = 6'ha == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1056; // @[Reg.scala 27:20]
  wire  _T_165 = 6'h9 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_995; // @[Reg.scala 27:20]
  wire  _T_163 = 6'h8 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_934; // @[Reg.scala 27:20]
  wire  _T_161 = 6'h7 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_873; // @[Reg.scala 27:20]
  wire  _T_159 = 6'h6 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_812; // @[Reg.scala 27:20]
  wire  _T_157 = 6'h5 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_751; // @[Reg.scala 27:20]
  wire  _T_155 = 6'h4 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_690; // @[Reg.scala 27:20]
  wire  _T_153 = 6'h3 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_629; // @[Reg.scala 27:20]
  wire  _T_151 = 6'h2 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_568; // @[Reg.scala 27:20]
  wire  _T_149 = 6'h1 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_507; // @[Reg.scala 27:20]
  reg  _T_446; // @[Reg.scala 27:20]
  wire  _T_150_0 = _T_149 ? _T_507 : _T_446; // @[Mux.scala 80:57]
  wire  _T_152_0 = _T_151 ? _T_568 : _T_150_0; // @[Mux.scala 80:57]
  wire  _T_154_0 = _T_153 ? _T_629 : _T_152_0; // @[Mux.scala 80:57]
  wire  _T_156_0 = _T_155 ? _T_690 : _T_154_0; // @[Mux.scala 80:57]
  wire  _T_158_0 = _T_157 ? _T_751 : _T_156_0; // @[Mux.scala 80:57]
  wire  _T_160_0 = _T_159 ? _T_812 : _T_158_0; // @[Mux.scala 80:57]
  wire  _T_162_0 = _T_161 ? _T_873 : _T_160_0; // @[Mux.scala 80:57]
  wire  _T_164_0 = _T_163 ? _T_934 : _T_162_0; // @[Mux.scala 80:57]
  wire  _T_166_0 = _T_165 ? _T_995 : _T_164_0; // @[Mux.scala 80:57]
  wire  _T_168_0 = _T_167 ? _T_1056 : _T_166_0; // @[Mux.scala 80:57]
  wire  _T_170_0 = _T_169 ? _T_1117 : _T_168_0; // @[Mux.scala 80:57]
  wire  _T_172_0 = _T_171 ? _T_1178 : _T_170_0; // @[Mux.scala 80:57]
  wire  _T_174_0 = _T_173 ? _T_1239 : _T_172_0; // @[Mux.scala 80:57]
  wire  _T_176_0 = _T_175 ? _T_1300 : _T_174_0; // @[Mux.scala 80:57]
  wire  _T_178_0 = _T_177 ? _T_1361 : _T_176_0; // @[Mux.scala 80:57]
  wire  _T_180_0 = _T_179 ? _T_1422 : _T_178_0; // @[Mux.scala 80:57]
  wire  _T_182_0 = _T_181 ? _T_1483 : _T_180_0; // @[Mux.scala 80:57]
  wire  _T_184_0 = _T_183 ? _T_1544 : _T_182_0; // @[Mux.scala 80:57]
  wire  _T_186_0 = _T_185 ? _T_1605 : _T_184_0; // @[Mux.scala 80:57]
  wire  _T_188_0 = _T_187 ? _T_1666 : _T_186_0; // @[Mux.scala 80:57]
  wire  _T_190_0 = _T_189 ? _T_1727 : _T_188_0; // @[Mux.scala 80:57]
  wire  _T_192_0 = _T_191 ? _T_1788 : _T_190_0; // @[Mux.scala 80:57]
  wire  _T_194_0 = _T_193 ? _T_1849 : _T_192_0; // @[Mux.scala 80:57]
  wire  _T_196_0 = _T_195 ? _T_1910 : _T_194_0; // @[Mux.scala 80:57]
  wire  _T_198_0 = _T_197 ? _T_1971 : _T_196_0; // @[Mux.scala 80:57]
  wire  _T_200_0 = _T_199 ? _T_2032 : _T_198_0; // @[Mux.scala 80:57]
  wire  _T_202_0 = _T_201 ? _T_2093 : _T_200_0; // @[Mux.scala 80:57]
  wire  _T_204_0 = _T_203 ? _T_2154 : _T_202_0; // @[Mux.scala 80:57]
  wire  _T_206_0 = _T_205 ? _T_2215 : _T_204_0; // @[Mux.scala 80:57]
  wire  _T_208_0 = _T_207 ? _T_2276 : _T_206_0; // @[Mux.scala 80:57]
  wire  _T_210_0 = _T_209 ? _T_2337 : _T_208_0; // @[Mux.scala 80:57]
  wire  _T_212_0 = _T_211 ? _T_2398 : _T_210_0; // @[Mux.scala 80:57]
  wire  _T_214_0 = _T_213 ? _T_2459 : _T_212_0; // @[Mux.scala 80:57]
  wire  _T_216_0 = _T_215 ? _T_2520 : _T_214_0; // @[Mux.scala 80:57]
  wire  _T_218_0 = _T_217 ? _T_2581 : _T_216_0; // @[Mux.scala 80:57]
  wire  _T_220_0 = _T_219 ? _T_2642 : _T_218_0; // @[Mux.scala 80:57]
  wire  _T_222_0 = _T_221 ? _T_2703 : _T_220_0; // @[Mux.scala 80:57]
  wire  _T_224_0 = _T_223 ? _T_2764 : _T_222_0; // @[Mux.scala 80:57]
  wire  _T_226_0 = _T_225 ? _T_2825 : _T_224_0; // @[Mux.scala 80:57]
  wire  _T_228_0 = _T_227 ? _T_2886 : _T_226_0; // @[Mux.scala 80:57]
  wire  _T_230_0 = _T_229 ? _T_2947 : _T_228_0; // @[Mux.scala 80:57]
  wire  _T_232_0 = _T_231 ? _T_3008 : _T_230_0; // @[Mux.scala 80:57]
  wire  _T_234_0 = _T_233 ? _T_3069 : _T_232_0; // @[Mux.scala 80:57]
  wire  _T_236_0 = _T_235 ? _T_3130 : _T_234_0; // @[Mux.scala 80:57]
  wire  _T_238_0 = _T_237 ? _T_3191 : _T_236_0; // @[Mux.scala 80:57]
  wire  _T_240_0 = _T_239 ? _T_3252 : _T_238_0; // @[Mux.scala 80:57]
  wire  _T_242_0 = _T_241 ? _T_3313 : _T_240_0; // @[Mux.scala 80:57]
  wire  _T_244_0 = _T_243 ? _T_3374 : _T_242_0; // @[Mux.scala 80:57]
  wire  _T_246_0 = _T_245 ? _T_3435 : _T_244_0; // @[Mux.scala 80:57]
  wire  _T_248_0 = _T_247 ? _T_3496 : _T_246_0; // @[Mux.scala 80:57]
  wire  _T_250_0 = _T_249 ? _T_3557 : _T_248_0; // @[Mux.scala 80:57]
  wire  _T_252_0 = _T_251 ? _T_3618 : _T_250_0; // @[Mux.scala 80:57]
  wire  _T_254_0 = _T_253 ? _T_3679 : _T_252_0; // @[Mux.scala 80:57]
  wire  _T_256_0 = _T_255 ? _T_3740 : _T_254_0; // @[Mux.scala 80:57]
  wire  _T_258_0 = _T_257 ? _T_3801 : _T_256_0; // @[Mux.scala 80:57]
  wire  _T_260_0 = _T_259 ? _T_3862 : _T_258_0; // @[Mux.scala 80:57]
  wire  _T_262_0 = _T_261 ? _T_3923 : _T_260_0; // @[Mux.scala 80:57]
  wire  _T_264_0 = _T_263 ? _T_3984 : _T_262_0; // @[Mux.scala 80:57]
  wire  _T_266_0 = _T_265 ? _T_4045 : _T_264_0; // @[Mux.scala 80:57]
  wire  _T_268_0 = _T_267 ? _T_4106 : _T_266_0; // @[Mux.scala 80:57]
  wire  _T_270_0 = _T_269 ? _T_4167 : _T_268_0; // @[Mux.scala 80:57]
  wire  _T_272_0 = _T_271 ? _T_4228 : _T_270_0; // @[Mux.scala 80:57]
  wire  _T_274_0 = _T_273 ? _T_4289 : _T_272_0; // @[Mux.scala 80:57]
  reg [21:0] _T_4281; // @[Reg.scala 27:20]
  reg [21:0] _T_4220; // @[Reg.scala 27:20]
  reg [21:0] _T_4159; // @[Reg.scala 27:20]
  reg [21:0] _T_4098; // @[Reg.scala 27:20]
  reg [21:0] _T_4037; // @[Reg.scala 27:20]
  reg [21:0] _T_3976; // @[Reg.scala 27:20]
  reg [21:0] _T_3915; // @[Reg.scala 27:20]
  reg [21:0] _T_3854; // @[Reg.scala 27:20]
  reg [21:0] _T_3793; // @[Reg.scala 27:20]
  reg [21:0] _T_3732; // @[Reg.scala 27:20]
  reg [21:0] _T_3671; // @[Reg.scala 27:20]
  reg [21:0] _T_3610; // @[Reg.scala 27:20]
  reg [21:0] _T_3549; // @[Reg.scala 27:20]
  reg [21:0] _T_3488; // @[Reg.scala 27:20]
  reg [21:0] _T_3427; // @[Reg.scala 27:20]
  reg [21:0] _T_3366; // @[Reg.scala 27:20]
  reg [21:0] _T_3305; // @[Reg.scala 27:20]
  reg [21:0] _T_3244; // @[Reg.scala 27:20]
  reg [21:0] _T_3183; // @[Reg.scala 27:20]
  reg [21:0] _T_3122; // @[Reg.scala 27:20]
  reg [21:0] _T_3061; // @[Reg.scala 27:20]
  reg [21:0] _T_3000; // @[Reg.scala 27:20]
  reg [21:0] _T_2939; // @[Reg.scala 27:20]
  reg [21:0] _T_2878; // @[Reg.scala 27:20]
  reg [21:0] _T_2817; // @[Reg.scala 27:20]
  reg [21:0] _T_2756; // @[Reg.scala 27:20]
  reg [21:0] _T_2695; // @[Reg.scala 27:20]
  reg [21:0] _T_2634; // @[Reg.scala 27:20]
  reg [21:0] _T_2573; // @[Reg.scala 27:20]
  reg [21:0] _T_2512; // @[Reg.scala 27:20]
  reg [21:0] _T_2451; // @[Reg.scala 27:20]
  reg [21:0] _T_2390; // @[Reg.scala 27:20]
  reg [21:0] _T_2329; // @[Reg.scala 27:20]
  reg [21:0] _T_2268; // @[Reg.scala 27:20]
  reg [21:0] _T_2207; // @[Reg.scala 27:20]
  reg [21:0] _T_2146; // @[Reg.scala 27:20]
  reg [21:0] _T_2085; // @[Reg.scala 27:20]
  reg [21:0] _T_2024; // @[Reg.scala 27:20]
  reg [21:0] _T_1963; // @[Reg.scala 27:20]
  reg [21:0] _T_1902; // @[Reg.scala 27:20]
  reg [21:0] _T_1841; // @[Reg.scala 27:20]
  reg [21:0] _T_1780; // @[Reg.scala 27:20]
  reg [21:0] _T_1719; // @[Reg.scala 27:20]
  reg [21:0] _T_1658; // @[Reg.scala 27:20]
  reg [21:0] _T_1597; // @[Reg.scala 27:20]
  reg [21:0] _T_1536; // @[Reg.scala 27:20]
  reg [21:0] _T_1475; // @[Reg.scala 27:20]
  reg [21:0] _T_1414; // @[Reg.scala 27:20]
  reg [21:0] _T_1353; // @[Reg.scala 27:20]
  reg [21:0] _T_1292; // @[Reg.scala 27:20]
  reg [21:0] _T_1231; // @[Reg.scala 27:20]
  reg [21:0] _T_1170; // @[Reg.scala 27:20]
  reg [21:0] _T_1109; // @[Reg.scala 27:20]
  reg [21:0] _T_1048; // @[Reg.scala 27:20]
  reg [21:0] _T_987; // @[Reg.scala 27:20]
  reg [21:0] _T_926; // @[Reg.scala 27:20]
  reg [21:0] _T_865; // @[Reg.scala 27:20]
  reg [21:0] _T_804; // @[Reg.scala 27:20]
  reg [21:0] _T_743; // @[Reg.scala 27:20]
  reg [21:0] _T_682; // @[Reg.scala 27:20]
  reg [21:0] _T_621; // @[Reg.scala 27:20]
  reg [21:0] _T_560; // @[Reg.scala 27:20]
  reg [21:0] _T_499; // @[Reg.scala 27:20]
  reg [21:0] _T_438; // @[Reg.scala 27:20]
  wire [21:0] _T_24_0 = _T_149 ? _T_499 : _T_438; // @[Mux.scala 80:57]
  wire [21:0] _T_26_0 = _T_151 ? _T_560 : _T_24_0; // @[Mux.scala 80:57]
  wire [21:0] _T_28_0 = _T_153 ? _T_621 : _T_26_0; // @[Mux.scala 80:57]
  wire [21:0] _T_30_0 = _T_155 ? _T_682 : _T_28_0; // @[Mux.scala 80:57]
  wire [21:0] _T_32_0 = _T_157 ? _T_743 : _T_30_0; // @[Mux.scala 80:57]
  wire [21:0] _T_34_0 = _T_159 ? _T_804 : _T_32_0; // @[Mux.scala 80:57]
  wire [21:0] _T_36_0 = _T_161 ? _T_865 : _T_34_0; // @[Mux.scala 80:57]
  wire [21:0] _T_38_0 = _T_163 ? _T_926 : _T_36_0; // @[Mux.scala 80:57]
  wire [21:0] _T_40_0 = _T_165 ? _T_987 : _T_38_0; // @[Mux.scala 80:57]
  wire [21:0] _T_42_0 = _T_167 ? _T_1048 : _T_40_0; // @[Mux.scala 80:57]
  wire [21:0] _T_44_0 = _T_169 ? _T_1109 : _T_42_0; // @[Mux.scala 80:57]
  wire [21:0] _T_46_0 = _T_171 ? _T_1170 : _T_44_0; // @[Mux.scala 80:57]
  wire [21:0] _T_48_0 = _T_173 ? _T_1231 : _T_46_0; // @[Mux.scala 80:57]
  wire [21:0] _T_50_0 = _T_175 ? _T_1292 : _T_48_0; // @[Mux.scala 80:57]
  wire [21:0] _T_52_0 = _T_177 ? _T_1353 : _T_50_0; // @[Mux.scala 80:57]
  wire [21:0] _T_54_0 = _T_179 ? _T_1414 : _T_52_0; // @[Mux.scala 80:57]
  wire [21:0] _T_56_0 = _T_181 ? _T_1475 : _T_54_0; // @[Mux.scala 80:57]
  wire [21:0] _T_58_0 = _T_183 ? _T_1536 : _T_56_0; // @[Mux.scala 80:57]
  wire [21:0] _T_60_0 = _T_185 ? _T_1597 : _T_58_0; // @[Mux.scala 80:57]
  wire [21:0] _T_62_0 = _T_187 ? _T_1658 : _T_60_0; // @[Mux.scala 80:57]
  wire [21:0] _T_64_0 = _T_189 ? _T_1719 : _T_62_0; // @[Mux.scala 80:57]
  wire [21:0] _T_66_0 = _T_191 ? _T_1780 : _T_64_0; // @[Mux.scala 80:57]
  wire [21:0] _T_68_0 = _T_193 ? _T_1841 : _T_66_0; // @[Mux.scala 80:57]
  wire [21:0] _T_70_0 = _T_195 ? _T_1902 : _T_68_0; // @[Mux.scala 80:57]
  wire [21:0] _T_72_0 = _T_197 ? _T_1963 : _T_70_0; // @[Mux.scala 80:57]
  wire [21:0] _T_74_0 = _T_199 ? _T_2024 : _T_72_0; // @[Mux.scala 80:57]
  wire [21:0] _T_76_0 = _T_201 ? _T_2085 : _T_74_0; // @[Mux.scala 80:57]
  wire [21:0] _T_78_0 = _T_203 ? _T_2146 : _T_76_0; // @[Mux.scala 80:57]
  wire [21:0] _T_80_0 = _T_205 ? _T_2207 : _T_78_0; // @[Mux.scala 80:57]
  wire [21:0] _T_82_0 = _T_207 ? _T_2268 : _T_80_0; // @[Mux.scala 80:57]
  wire [21:0] _T_84_0 = _T_209 ? _T_2329 : _T_82_0; // @[Mux.scala 80:57]
  wire [21:0] _T_86_0 = _T_211 ? _T_2390 : _T_84_0; // @[Mux.scala 80:57]
  wire [21:0] _T_88_0 = _T_213 ? _T_2451 : _T_86_0; // @[Mux.scala 80:57]
  wire [21:0] _T_90_0 = _T_215 ? _T_2512 : _T_88_0; // @[Mux.scala 80:57]
  wire [21:0] _T_92_0 = _T_217 ? _T_2573 : _T_90_0; // @[Mux.scala 80:57]
  wire [21:0] _T_94_0 = _T_219 ? _T_2634 : _T_92_0; // @[Mux.scala 80:57]
  wire [21:0] _T_96_0 = _T_221 ? _T_2695 : _T_94_0; // @[Mux.scala 80:57]
  wire [21:0] _T_98_0 = _T_223 ? _T_2756 : _T_96_0; // @[Mux.scala 80:57]
  wire [21:0] _T_100_0 = _T_225 ? _T_2817 : _T_98_0; // @[Mux.scala 80:57]
  wire [21:0] _T_102_0 = _T_227 ? _T_2878 : _T_100_0; // @[Mux.scala 80:57]
  wire [21:0] _T_104_0 = _T_229 ? _T_2939 : _T_102_0; // @[Mux.scala 80:57]
  wire [21:0] _T_106_0 = _T_231 ? _T_3000 : _T_104_0; // @[Mux.scala 80:57]
  wire [21:0] _T_108_0 = _T_233 ? _T_3061 : _T_106_0; // @[Mux.scala 80:57]
  wire [21:0] _T_110_0 = _T_235 ? _T_3122 : _T_108_0; // @[Mux.scala 80:57]
  wire [21:0] _T_112_0 = _T_237 ? _T_3183 : _T_110_0; // @[Mux.scala 80:57]
  wire [21:0] _T_114_0 = _T_239 ? _T_3244 : _T_112_0; // @[Mux.scala 80:57]
  wire [21:0] _T_116_0 = _T_241 ? _T_3305 : _T_114_0; // @[Mux.scala 80:57]
  wire [21:0] _T_118_0 = _T_243 ? _T_3366 : _T_116_0; // @[Mux.scala 80:57]
  wire [21:0] _T_120_0 = _T_245 ? _T_3427 : _T_118_0; // @[Mux.scala 80:57]
  wire [21:0] _T_122_0 = _T_247 ? _T_3488 : _T_120_0; // @[Mux.scala 80:57]
  wire [21:0] _T_124_0 = _T_249 ? _T_3549 : _T_122_0; // @[Mux.scala 80:57]
  wire [21:0] _T_126_0 = _T_251 ? _T_3610 : _T_124_0; // @[Mux.scala 80:57]
  wire [21:0] _T_128_0 = _T_253 ? _T_3671 : _T_126_0; // @[Mux.scala 80:57]
  wire [21:0] _T_130_0 = _T_255 ? _T_3732 : _T_128_0; // @[Mux.scala 80:57]
  wire [21:0] _T_132_0 = _T_257 ? _T_3793 : _T_130_0; // @[Mux.scala 80:57]
  wire [21:0] _T_134_0 = _T_259 ? _T_3854 : _T_132_0; // @[Mux.scala 80:57]
  wire [21:0] _T_136_0 = _T_261 ? _T_3915 : _T_134_0; // @[Mux.scala 80:57]
  wire [21:0] _T_138_0 = _T_263 ? _T_3976 : _T_136_0; // @[Mux.scala 80:57]
  wire [21:0] _T_140_0 = _T_265 ? _T_4037 : _T_138_0; // @[Mux.scala 80:57]
  wire [21:0] _T_142_0 = _T_267 ? _T_4098 : _T_140_0; // @[Mux.scala 80:57]
  wire [21:0] _T_144_0 = _T_269 ? _T_4159 : _T_142_0; // @[Mux.scala 80:57]
  wire [21:0] _T_146_0 = _T_271 ? _T_4220 : _T_144_0; // @[Mux.scala 80:57]
  wire [21:0] _T_148_0 = _T_273 ? _T_4281 : _T_146_0; // @[Mux.scala 80:57]
  wire  _T_275 = _T_148_0 == io_cacheIn_addr[31:10]; // @[Cache.scala 446:76]
  wire  _T_276 = _T_274_0 & _T_275; // @[Cache.scala 446:60]
  reg  _T_4303; // @[Reg.scala 27:20]
  reg  _T_4242; // @[Reg.scala 27:20]
  reg  _T_4181; // @[Reg.scala 27:20]
  reg  _T_4120; // @[Reg.scala 27:20]
  reg  _T_4059; // @[Reg.scala 27:20]
  reg  _T_3998; // @[Reg.scala 27:20]
  reg  _T_3937; // @[Reg.scala 27:20]
  reg  _T_3876; // @[Reg.scala 27:20]
  reg  _T_3815; // @[Reg.scala 27:20]
  reg  _T_3754; // @[Reg.scala 27:20]
  reg  _T_3693; // @[Reg.scala 27:20]
  reg  _T_3632; // @[Reg.scala 27:20]
  reg  _T_3571; // @[Reg.scala 27:20]
  reg  _T_3510; // @[Reg.scala 27:20]
  reg  _T_3449; // @[Reg.scala 27:20]
  reg  _T_3388; // @[Reg.scala 27:20]
  reg  _T_3327; // @[Reg.scala 27:20]
  reg  _T_3266; // @[Reg.scala 27:20]
  reg  _T_3205; // @[Reg.scala 27:20]
  reg  _T_3144; // @[Reg.scala 27:20]
  reg  _T_3083; // @[Reg.scala 27:20]
  reg  _T_3022; // @[Reg.scala 27:20]
  reg  _T_2961; // @[Reg.scala 27:20]
  reg  _T_2900; // @[Reg.scala 27:20]
  reg  _T_2839; // @[Reg.scala 27:20]
  reg  _T_2778; // @[Reg.scala 27:20]
  reg  _T_2717; // @[Reg.scala 27:20]
  reg  _T_2656; // @[Reg.scala 27:20]
  reg  _T_2595; // @[Reg.scala 27:20]
  reg  _T_2534; // @[Reg.scala 27:20]
  reg  _T_2473; // @[Reg.scala 27:20]
  reg  _T_2412; // @[Reg.scala 27:20]
  reg  _T_2351; // @[Reg.scala 27:20]
  reg  _T_2290; // @[Reg.scala 27:20]
  reg  _T_2229; // @[Reg.scala 27:20]
  reg  _T_2168; // @[Reg.scala 27:20]
  reg  _T_2107; // @[Reg.scala 27:20]
  reg  _T_2046; // @[Reg.scala 27:20]
  reg  _T_1985; // @[Reg.scala 27:20]
  reg  _T_1924; // @[Reg.scala 27:20]
  reg  _T_1863; // @[Reg.scala 27:20]
  reg  _T_1802; // @[Reg.scala 27:20]
  reg  _T_1741; // @[Reg.scala 27:20]
  reg  _T_1680; // @[Reg.scala 27:20]
  reg  _T_1619; // @[Reg.scala 27:20]
  reg  _T_1558; // @[Reg.scala 27:20]
  reg  _T_1497; // @[Reg.scala 27:20]
  reg  _T_1436; // @[Reg.scala 27:20]
  reg  _T_1375; // @[Reg.scala 27:20]
  reg  _T_1314; // @[Reg.scala 27:20]
  reg  _T_1253; // @[Reg.scala 27:20]
  reg  _T_1192; // @[Reg.scala 27:20]
  reg  _T_1131; // @[Reg.scala 27:20]
  reg  _T_1070; // @[Reg.scala 27:20]
  reg  _T_1009; // @[Reg.scala 27:20]
  reg  _T_948; // @[Reg.scala 27:20]
  reg  _T_887; // @[Reg.scala 27:20]
  reg  _T_826; // @[Reg.scala 27:20]
  reg  _T_765; // @[Reg.scala 27:20]
  reg  _T_704; // @[Reg.scala 27:20]
  reg  _T_643; // @[Reg.scala 27:20]
  reg  _T_582; // @[Reg.scala 27:20]
  reg  _T_521; // @[Reg.scala 27:20]
  reg  _T_460; // @[Reg.scala 27:20]
  wire  _T_150_1 = _T_149 ? _T_521 : _T_460; // @[Mux.scala 80:57]
  wire  _T_152_1 = _T_151 ? _T_582 : _T_150_1; // @[Mux.scala 80:57]
  wire  _T_154_1 = _T_153 ? _T_643 : _T_152_1; // @[Mux.scala 80:57]
  wire  _T_156_1 = _T_155 ? _T_704 : _T_154_1; // @[Mux.scala 80:57]
  wire  _T_158_1 = _T_157 ? _T_765 : _T_156_1; // @[Mux.scala 80:57]
  wire  _T_160_1 = _T_159 ? _T_826 : _T_158_1; // @[Mux.scala 80:57]
  wire  _T_162_1 = _T_161 ? _T_887 : _T_160_1; // @[Mux.scala 80:57]
  wire  _T_164_1 = _T_163 ? _T_948 : _T_162_1; // @[Mux.scala 80:57]
  wire  _T_166_1 = _T_165 ? _T_1009 : _T_164_1; // @[Mux.scala 80:57]
  wire  _T_168_1 = _T_167 ? _T_1070 : _T_166_1; // @[Mux.scala 80:57]
  wire  _T_170_1 = _T_169 ? _T_1131 : _T_168_1; // @[Mux.scala 80:57]
  wire  _T_172_1 = _T_171 ? _T_1192 : _T_170_1; // @[Mux.scala 80:57]
  wire  _T_174_1 = _T_173 ? _T_1253 : _T_172_1; // @[Mux.scala 80:57]
  wire  _T_176_1 = _T_175 ? _T_1314 : _T_174_1; // @[Mux.scala 80:57]
  wire  _T_178_1 = _T_177 ? _T_1375 : _T_176_1; // @[Mux.scala 80:57]
  wire  _T_180_1 = _T_179 ? _T_1436 : _T_178_1; // @[Mux.scala 80:57]
  wire  _T_182_1 = _T_181 ? _T_1497 : _T_180_1; // @[Mux.scala 80:57]
  wire  _T_184_1 = _T_183 ? _T_1558 : _T_182_1; // @[Mux.scala 80:57]
  wire  _T_186_1 = _T_185 ? _T_1619 : _T_184_1; // @[Mux.scala 80:57]
  wire  _T_188_1 = _T_187 ? _T_1680 : _T_186_1; // @[Mux.scala 80:57]
  wire  _T_190_1 = _T_189 ? _T_1741 : _T_188_1; // @[Mux.scala 80:57]
  wire  _T_192_1 = _T_191 ? _T_1802 : _T_190_1; // @[Mux.scala 80:57]
  wire  _T_194_1 = _T_193 ? _T_1863 : _T_192_1; // @[Mux.scala 80:57]
  wire  _T_196_1 = _T_195 ? _T_1924 : _T_194_1; // @[Mux.scala 80:57]
  wire  _T_198_1 = _T_197 ? _T_1985 : _T_196_1; // @[Mux.scala 80:57]
  wire  _T_200_1 = _T_199 ? _T_2046 : _T_198_1; // @[Mux.scala 80:57]
  wire  _T_202_1 = _T_201 ? _T_2107 : _T_200_1; // @[Mux.scala 80:57]
  wire  _T_204_1 = _T_203 ? _T_2168 : _T_202_1; // @[Mux.scala 80:57]
  wire  _T_206_1 = _T_205 ? _T_2229 : _T_204_1; // @[Mux.scala 80:57]
  wire  _T_208_1 = _T_207 ? _T_2290 : _T_206_1; // @[Mux.scala 80:57]
  wire  _T_210_1 = _T_209 ? _T_2351 : _T_208_1; // @[Mux.scala 80:57]
  wire  _T_212_1 = _T_211 ? _T_2412 : _T_210_1; // @[Mux.scala 80:57]
  wire  _T_214_1 = _T_213 ? _T_2473 : _T_212_1; // @[Mux.scala 80:57]
  wire  _T_216_1 = _T_215 ? _T_2534 : _T_214_1; // @[Mux.scala 80:57]
  wire  _T_218_1 = _T_217 ? _T_2595 : _T_216_1; // @[Mux.scala 80:57]
  wire  _T_220_1 = _T_219 ? _T_2656 : _T_218_1; // @[Mux.scala 80:57]
  wire  _T_222_1 = _T_221 ? _T_2717 : _T_220_1; // @[Mux.scala 80:57]
  wire  _T_224_1 = _T_223 ? _T_2778 : _T_222_1; // @[Mux.scala 80:57]
  wire  _T_226_1 = _T_225 ? _T_2839 : _T_224_1; // @[Mux.scala 80:57]
  wire  _T_228_1 = _T_227 ? _T_2900 : _T_226_1; // @[Mux.scala 80:57]
  wire  _T_230_1 = _T_229 ? _T_2961 : _T_228_1; // @[Mux.scala 80:57]
  wire  _T_232_1 = _T_231 ? _T_3022 : _T_230_1; // @[Mux.scala 80:57]
  wire  _T_234_1 = _T_233 ? _T_3083 : _T_232_1; // @[Mux.scala 80:57]
  wire  _T_236_1 = _T_235 ? _T_3144 : _T_234_1; // @[Mux.scala 80:57]
  wire  _T_238_1 = _T_237 ? _T_3205 : _T_236_1; // @[Mux.scala 80:57]
  wire  _T_240_1 = _T_239 ? _T_3266 : _T_238_1; // @[Mux.scala 80:57]
  wire  _T_242_1 = _T_241 ? _T_3327 : _T_240_1; // @[Mux.scala 80:57]
  wire  _T_244_1 = _T_243 ? _T_3388 : _T_242_1; // @[Mux.scala 80:57]
  wire  _T_246_1 = _T_245 ? _T_3449 : _T_244_1; // @[Mux.scala 80:57]
  wire  _T_248_1 = _T_247 ? _T_3510 : _T_246_1; // @[Mux.scala 80:57]
  wire  _T_250_1 = _T_249 ? _T_3571 : _T_248_1; // @[Mux.scala 80:57]
  wire  _T_252_1 = _T_251 ? _T_3632 : _T_250_1; // @[Mux.scala 80:57]
  wire  _T_254_1 = _T_253 ? _T_3693 : _T_252_1; // @[Mux.scala 80:57]
  wire  _T_256_1 = _T_255 ? _T_3754 : _T_254_1; // @[Mux.scala 80:57]
  wire  _T_258_1 = _T_257 ? _T_3815 : _T_256_1; // @[Mux.scala 80:57]
  wire  _T_260_1 = _T_259 ? _T_3876 : _T_258_1; // @[Mux.scala 80:57]
  wire  _T_262_1 = _T_261 ? _T_3937 : _T_260_1; // @[Mux.scala 80:57]
  wire  _T_264_1 = _T_263 ? _T_3998 : _T_262_1; // @[Mux.scala 80:57]
  wire  _T_266_1 = _T_265 ? _T_4059 : _T_264_1; // @[Mux.scala 80:57]
  wire  _T_268_1 = _T_267 ? _T_4120 : _T_266_1; // @[Mux.scala 80:57]
  wire  _T_270_1 = _T_269 ? _T_4181 : _T_268_1; // @[Mux.scala 80:57]
  wire  _T_272_1 = _T_271 ? _T_4242 : _T_270_1; // @[Mux.scala 80:57]
  wire  _T_274_1 = _T_273 ? _T_4303 : _T_272_1; // @[Mux.scala 80:57]
  reg [21:0] _T_4295; // @[Reg.scala 27:20]
  reg [21:0] _T_4234; // @[Reg.scala 27:20]
  reg [21:0] _T_4173; // @[Reg.scala 27:20]
  reg [21:0] _T_4112; // @[Reg.scala 27:20]
  reg [21:0] _T_4051; // @[Reg.scala 27:20]
  reg [21:0] _T_3990; // @[Reg.scala 27:20]
  reg [21:0] _T_3929; // @[Reg.scala 27:20]
  reg [21:0] _T_3868; // @[Reg.scala 27:20]
  reg [21:0] _T_3807; // @[Reg.scala 27:20]
  reg [21:0] _T_3746; // @[Reg.scala 27:20]
  reg [21:0] _T_3685; // @[Reg.scala 27:20]
  reg [21:0] _T_3624; // @[Reg.scala 27:20]
  reg [21:0] _T_3563; // @[Reg.scala 27:20]
  reg [21:0] _T_3502; // @[Reg.scala 27:20]
  reg [21:0] _T_3441; // @[Reg.scala 27:20]
  reg [21:0] _T_3380; // @[Reg.scala 27:20]
  reg [21:0] _T_3319; // @[Reg.scala 27:20]
  reg [21:0] _T_3258; // @[Reg.scala 27:20]
  reg [21:0] _T_3197; // @[Reg.scala 27:20]
  reg [21:0] _T_3136; // @[Reg.scala 27:20]
  reg [21:0] _T_3075; // @[Reg.scala 27:20]
  reg [21:0] _T_3014; // @[Reg.scala 27:20]
  reg [21:0] _T_2953; // @[Reg.scala 27:20]
  reg [21:0] _T_2892; // @[Reg.scala 27:20]
  reg [21:0] _T_2831; // @[Reg.scala 27:20]
  reg [21:0] _T_2770; // @[Reg.scala 27:20]
  reg [21:0] _T_2709; // @[Reg.scala 27:20]
  reg [21:0] _T_2648; // @[Reg.scala 27:20]
  reg [21:0] _T_2587; // @[Reg.scala 27:20]
  reg [21:0] _T_2526; // @[Reg.scala 27:20]
  reg [21:0] _T_2465; // @[Reg.scala 27:20]
  reg [21:0] _T_2404; // @[Reg.scala 27:20]
  reg [21:0] _T_2343; // @[Reg.scala 27:20]
  reg [21:0] _T_2282; // @[Reg.scala 27:20]
  reg [21:0] _T_2221; // @[Reg.scala 27:20]
  reg [21:0] _T_2160; // @[Reg.scala 27:20]
  reg [21:0] _T_2099; // @[Reg.scala 27:20]
  reg [21:0] _T_2038; // @[Reg.scala 27:20]
  reg [21:0] _T_1977; // @[Reg.scala 27:20]
  reg [21:0] _T_1916; // @[Reg.scala 27:20]
  reg [21:0] _T_1855; // @[Reg.scala 27:20]
  reg [21:0] _T_1794; // @[Reg.scala 27:20]
  reg [21:0] _T_1733; // @[Reg.scala 27:20]
  reg [21:0] _T_1672; // @[Reg.scala 27:20]
  reg [21:0] _T_1611; // @[Reg.scala 27:20]
  reg [21:0] _T_1550; // @[Reg.scala 27:20]
  reg [21:0] _T_1489; // @[Reg.scala 27:20]
  reg [21:0] _T_1428; // @[Reg.scala 27:20]
  reg [21:0] _T_1367; // @[Reg.scala 27:20]
  reg [21:0] _T_1306; // @[Reg.scala 27:20]
  reg [21:0] _T_1245; // @[Reg.scala 27:20]
  reg [21:0] _T_1184; // @[Reg.scala 27:20]
  reg [21:0] _T_1123; // @[Reg.scala 27:20]
  reg [21:0] _T_1062; // @[Reg.scala 27:20]
  reg [21:0] _T_1001; // @[Reg.scala 27:20]
  reg [21:0] _T_940; // @[Reg.scala 27:20]
  reg [21:0] _T_879; // @[Reg.scala 27:20]
  reg [21:0] _T_818; // @[Reg.scala 27:20]
  reg [21:0] _T_757; // @[Reg.scala 27:20]
  reg [21:0] _T_696; // @[Reg.scala 27:20]
  reg [21:0] _T_635; // @[Reg.scala 27:20]
  reg [21:0] _T_574; // @[Reg.scala 27:20]
  reg [21:0] _T_513; // @[Reg.scala 27:20]
  reg [21:0] _T_452; // @[Reg.scala 27:20]
  wire [21:0] _T_24_1 = _T_149 ? _T_513 : _T_452; // @[Mux.scala 80:57]
  wire [21:0] _T_26_1 = _T_151 ? _T_574 : _T_24_1; // @[Mux.scala 80:57]
  wire [21:0] _T_28_1 = _T_153 ? _T_635 : _T_26_1; // @[Mux.scala 80:57]
  wire [21:0] _T_30_1 = _T_155 ? _T_696 : _T_28_1; // @[Mux.scala 80:57]
  wire [21:0] _T_32_1 = _T_157 ? _T_757 : _T_30_1; // @[Mux.scala 80:57]
  wire [21:0] _T_34_1 = _T_159 ? _T_818 : _T_32_1; // @[Mux.scala 80:57]
  wire [21:0] _T_36_1 = _T_161 ? _T_879 : _T_34_1; // @[Mux.scala 80:57]
  wire [21:0] _T_38_1 = _T_163 ? _T_940 : _T_36_1; // @[Mux.scala 80:57]
  wire [21:0] _T_40_1 = _T_165 ? _T_1001 : _T_38_1; // @[Mux.scala 80:57]
  wire [21:0] _T_42_1 = _T_167 ? _T_1062 : _T_40_1; // @[Mux.scala 80:57]
  wire [21:0] _T_44_1 = _T_169 ? _T_1123 : _T_42_1; // @[Mux.scala 80:57]
  wire [21:0] _T_46_1 = _T_171 ? _T_1184 : _T_44_1; // @[Mux.scala 80:57]
  wire [21:0] _T_48_1 = _T_173 ? _T_1245 : _T_46_1; // @[Mux.scala 80:57]
  wire [21:0] _T_50_1 = _T_175 ? _T_1306 : _T_48_1; // @[Mux.scala 80:57]
  wire [21:0] _T_52_1 = _T_177 ? _T_1367 : _T_50_1; // @[Mux.scala 80:57]
  wire [21:0] _T_54_1 = _T_179 ? _T_1428 : _T_52_1; // @[Mux.scala 80:57]
  wire [21:0] _T_56_1 = _T_181 ? _T_1489 : _T_54_1; // @[Mux.scala 80:57]
  wire [21:0] _T_58_1 = _T_183 ? _T_1550 : _T_56_1; // @[Mux.scala 80:57]
  wire [21:0] _T_60_1 = _T_185 ? _T_1611 : _T_58_1; // @[Mux.scala 80:57]
  wire [21:0] _T_62_1 = _T_187 ? _T_1672 : _T_60_1; // @[Mux.scala 80:57]
  wire [21:0] _T_64_1 = _T_189 ? _T_1733 : _T_62_1; // @[Mux.scala 80:57]
  wire [21:0] _T_66_1 = _T_191 ? _T_1794 : _T_64_1; // @[Mux.scala 80:57]
  wire [21:0] _T_68_1 = _T_193 ? _T_1855 : _T_66_1; // @[Mux.scala 80:57]
  wire [21:0] _T_70_1 = _T_195 ? _T_1916 : _T_68_1; // @[Mux.scala 80:57]
  wire [21:0] _T_72_1 = _T_197 ? _T_1977 : _T_70_1; // @[Mux.scala 80:57]
  wire [21:0] _T_74_1 = _T_199 ? _T_2038 : _T_72_1; // @[Mux.scala 80:57]
  wire [21:0] _T_76_1 = _T_201 ? _T_2099 : _T_74_1; // @[Mux.scala 80:57]
  wire [21:0] _T_78_1 = _T_203 ? _T_2160 : _T_76_1; // @[Mux.scala 80:57]
  wire [21:0] _T_80_1 = _T_205 ? _T_2221 : _T_78_1; // @[Mux.scala 80:57]
  wire [21:0] _T_82_1 = _T_207 ? _T_2282 : _T_80_1; // @[Mux.scala 80:57]
  wire [21:0] _T_84_1 = _T_209 ? _T_2343 : _T_82_1; // @[Mux.scala 80:57]
  wire [21:0] _T_86_1 = _T_211 ? _T_2404 : _T_84_1; // @[Mux.scala 80:57]
  wire [21:0] _T_88_1 = _T_213 ? _T_2465 : _T_86_1; // @[Mux.scala 80:57]
  wire [21:0] _T_90_1 = _T_215 ? _T_2526 : _T_88_1; // @[Mux.scala 80:57]
  wire [21:0] _T_92_1 = _T_217 ? _T_2587 : _T_90_1; // @[Mux.scala 80:57]
  wire [21:0] _T_94_1 = _T_219 ? _T_2648 : _T_92_1; // @[Mux.scala 80:57]
  wire [21:0] _T_96_1 = _T_221 ? _T_2709 : _T_94_1; // @[Mux.scala 80:57]
  wire [21:0] _T_98_1 = _T_223 ? _T_2770 : _T_96_1; // @[Mux.scala 80:57]
  wire [21:0] _T_100_1 = _T_225 ? _T_2831 : _T_98_1; // @[Mux.scala 80:57]
  wire [21:0] _T_102_1 = _T_227 ? _T_2892 : _T_100_1; // @[Mux.scala 80:57]
  wire [21:0] _T_104_1 = _T_229 ? _T_2953 : _T_102_1; // @[Mux.scala 80:57]
  wire [21:0] _T_106_1 = _T_231 ? _T_3014 : _T_104_1; // @[Mux.scala 80:57]
  wire [21:0] _T_108_1 = _T_233 ? _T_3075 : _T_106_1; // @[Mux.scala 80:57]
  wire [21:0] _T_110_1 = _T_235 ? _T_3136 : _T_108_1; // @[Mux.scala 80:57]
  wire [21:0] _T_112_1 = _T_237 ? _T_3197 : _T_110_1; // @[Mux.scala 80:57]
  wire [21:0] _T_114_1 = _T_239 ? _T_3258 : _T_112_1; // @[Mux.scala 80:57]
  wire [21:0] _T_116_1 = _T_241 ? _T_3319 : _T_114_1; // @[Mux.scala 80:57]
  wire [21:0] _T_118_1 = _T_243 ? _T_3380 : _T_116_1; // @[Mux.scala 80:57]
  wire [21:0] _T_120_1 = _T_245 ? _T_3441 : _T_118_1; // @[Mux.scala 80:57]
  wire [21:0] _T_122_1 = _T_247 ? _T_3502 : _T_120_1; // @[Mux.scala 80:57]
  wire [21:0] _T_124_1 = _T_249 ? _T_3563 : _T_122_1; // @[Mux.scala 80:57]
  wire [21:0] _T_126_1 = _T_251 ? _T_3624 : _T_124_1; // @[Mux.scala 80:57]
  wire [21:0] _T_128_1 = _T_253 ? _T_3685 : _T_126_1; // @[Mux.scala 80:57]
  wire [21:0] _T_130_1 = _T_255 ? _T_3746 : _T_128_1; // @[Mux.scala 80:57]
  wire [21:0] _T_132_1 = _T_257 ? _T_3807 : _T_130_1; // @[Mux.scala 80:57]
  wire [21:0] _T_134_1 = _T_259 ? _T_3868 : _T_132_1; // @[Mux.scala 80:57]
  wire [21:0] _T_136_1 = _T_261 ? _T_3929 : _T_134_1; // @[Mux.scala 80:57]
  wire [21:0] _T_138_1 = _T_263 ? _T_3990 : _T_136_1; // @[Mux.scala 80:57]
  wire [21:0] _T_140_1 = _T_265 ? _T_4051 : _T_138_1; // @[Mux.scala 80:57]
  wire [21:0] _T_142_1 = _T_267 ? _T_4112 : _T_140_1; // @[Mux.scala 80:57]
  wire [21:0] _T_144_1 = _T_269 ? _T_4173 : _T_142_1; // @[Mux.scala 80:57]
  wire [21:0] _T_146_1 = _T_271 ? _T_4234 : _T_144_1; // @[Mux.scala 80:57]
  wire [21:0] _T_148_1 = _T_273 ? _T_4295 : _T_146_1; // @[Mux.scala 80:57]
  wire  _T_277 = _T_148_1 == io_cacheIn_addr[31:10]; // @[Cache.scala 446:76]
  wire  _T_278 = _T_274_1 & _T_277; // @[Cache.scala 446:60]
  wire  _T_284 = _T_276 | _T_278; // @[Cache.scala 447:49]
  reg  _T_4317; // @[Reg.scala 27:20]
  reg  _T_4256; // @[Reg.scala 27:20]
  reg  _T_4195; // @[Reg.scala 27:20]
  reg  _T_4134; // @[Reg.scala 27:20]
  reg  _T_4073; // @[Reg.scala 27:20]
  reg  _T_4012; // @[Reg.scala 27:20]
  reg  _T_3951; // @[Reg.scala 27:20]
  reg  _T_3890; // @[Reg.scala 27:20]
  reg  _T_3829; // @[Reg.scala 27:20]
  reg  _T_3768; // @[Reg.scala 27:20]
  reg  _T_3707; // @[Reg.scala 27:20]
  reg  _T_3646; // @[Reg.scala 27:20]
  reg  _T_3585; // @[Reg.scala 27:20]
  reg  _T_3524; // @[Reg.scala 27:20]
  reg  _T_3463; // @[Reg.scala 27:20]
  reg  _T_3402; // @[Reg.scala 27:20]
  reg  _T_3341; // @[Reg.scala 27:20]
  reg  _T_3280; // @[Reg.scala 27:20]
  reg  _T_3219; // @[Reg.scala 27:20]
  reg  _T_3158; // @[Reg.scala 27:20]
  reg  _T_3097; // @[Reg.scala 27:20]
  reg  _T_3036; // @[Reg.scala 27:20]
  reg  _T_2975; // @[Reg.scala 27:20]
  reg  _T_2914; // @[Reg.scala 27:20]
  reg  _T_2853; // @[Reg.scala 27:20]
  reg  _T_2792; // @[Reg.scala 27:20]
  reg  _T_2731; // @[Reg.scala 27:20]
  reg  _T_2670; // @[Reg.scala 27:20]
  reg  _T_2609; // @[Reg.scala 27:20]
  reg  _T_2548; // @[Reg.scala 27:20]
  reg  _T_2487; // @[Reg.scala 27:20]
  reg  _T_2426; // @[Reg.scala 27:20]
  reg  _T_2365; // @[Reg.scala 27:20]
  reg  _T_2304; // @[Reg.scala 27:20]
  reg  _T_2243; // @[Reg.scala 27:20]
  reg  _T_2182; // @[Reg.scala 27:20]
  reg  _T_2121; // @[Reg.scala 27:20]
  reg  _T_2060; // @[Reg.scala 27:20]
  reg  _T_1999; // @[Reg.scala 27:20]
  reg  _T_1938; // @[Reg.scala 27:20]
  reg  _T_1877; // @[Reg.scala 27:20]
  reg  _T_1816; // @[Reg.scala 27:20]
  reg  _T_1755; // @[Reg.scala 27:20]
  reg  _T_1694; // @[Reg.scala 27:20]
  reg  _T_1633; // @[Reg.scala 27:20]
  reg  _T_1572; // @[Reg.scala 27:20]
  reg  _T_1511; // @[Reg.scala 27:20]
  reg  _T_1450; // @[Reg.scala 27:20]
  reg  _T_1389; // @[Reg.scala 27:20]
  reg  _T_1328; // @[Reg.scala 27:20]
  reg  _T_1267; // @[Reg.scala 27:20]
  reg  _T_1206; // @[Reg.scala 27:20]
  reg  _T_1145; // @[Reg.scala 27:20]
  reg  _T_1084; // @[Reg.scala 27:20]
  reg  _T_1023; // @[Reg.scala 27:20]
  reg  _T_962; // @[Reg.scala 27:20]
  reg  _T_901; // @[Reg.scala 27:20]
  reg  _T_840; // @[Reg.scala 27:20]
  reg  _T_779; // @[Reg.scala 27:20]
  reg  _T_718; // @[Reg.scala 27:20]
  reg  _T_657; // @[Reg.scala 27:20]
  reg  _T_596; // @[Reg.scala 27:20]
  reg  _T_535; // @[Reg.scala 27:20]
  reg  _T_474; // @[Reg.scala 27:20]
  wire  _T_150_2 = _T_149 ? _T_535 : _T_474; // @[Mux.scala 80:57]
  wire  _T_152_2 = _T_151 ? _T_596 : _T_150_2; // @[Mux.scala 80:57]
  wire  _T_154_2 = _T_153 ? _T_657 : _T_152_2; // @[Mux.scala 80:57]
  wire  _T_156_2 = _T_155 ? _T_718 : _T_154_2; // @[Mux.scala 80:57]
  wire  _T_158_2 = _T_157 ? _T_779 : _T_156_2; // @[Mux.scala 80:57]
  wire  _T_160_2 = _T_159 ? _T_840 : _T_158_2; // @[Mux.scala 80:57]
  wire  _T_162_2 = _T_161 ? _T_901 : _T_160_2; // @[Mux.scala 80:57]
  wire  _T_164_2 = _T_163 ? _T_962 : _T_162_2; // @[Mux.scala 80:57]
  wire  _T_166_2 = _T_165 ? _T_1023 : _T_164_2; // @[Mux.scala 80:57]
  wire  _T_168_2 = _T_167 ? _T_1084 : _T_166_2; // @[Mux.scala 80:57]
  wire  _T_170_2 = _T_169 ? _T_1145 : _T_168_2; // @[Mux.scala 80:57]
  wire  _T_172_2 = _T_171 ? _T_1206 : _T_170_2; // @[Mux.scala 80:57]
  wire  _T_174_2 = _T_173 ? _T_1267 : _T_172_2; // @[Mux.scala 80:57]
  wire  _T_176_2 = _T_175 ? _T_1328 : _T_174_2; // @[Mux.scala 80:57]
  wire  _T_178_2 = _T_177 ? _T_1389 : _T_176_2; // @[Mux.scala 80:57]
  wire  _T_180_2 = _T_179 ? _T_1450 : _T_178_2; // @[Mux.scala 80:57]
  wire  _T_182_2 = _T_181 ? _T_1511 : _T_180_2; // @[Mux.scala 80:57]
  wire  _T_184_2 = _T_183 ? _T_1572 : _T_182_2; // @[Mux.scala 80:57]
  wire  _T_186_2 = _T_185 ? _T_1633 : _T_184_2; // @[Mux.scala 80:57]
  wire  _T_188_2 = _T_187 ? _T_1694 : _T_186_2; // @[Mux.scala 80:57]
  wire  _T_190_2 = _T_189 ? _T_1755 : _T_188_2; // @[Mux.scala 80:57]
  wire  _T_192_2 = _T_191 ? _T_1816 : _T_190_2; // @[Mux.scala 80:57]
  wire  _T_194_2 = _T_193 ? _T_1877 : _T_192_2; // @[Mux.scala 80:57]
  wire  _T_196_2 = _T_195 ? _T_1938 : _T_194_2; // @[Mux.scala 80:57]
  wire  _T_198_2 = _T_197 ? _T_1999 : _T_196_2; // @[Mux.scala 80:57]
  wire  _T_200_2 = _T_199 ? _T_2060 : _T_198_2; // @[Mux.scala 80:57]
  wire  _T_202_2 = _T_201 ? _T_2121 : _T_200_2; // @[Mux.scala 80:57]
  wire  _T_204_2 = _T_203 ? _T_2182 : _T_202_2; // @[Mux.scala 80:57]
  wire  _T_206_2 = _T_205 ? _T_2243 : _T_204_2; // @[Mux.scala 80:57]
  wire  _T_208_2 = _T_207 ? _T_2304 : _T_206_2; // @[Mux.scala 80:57]
  wire  _T_210_2 = _T_209 ? _T_2365 : _T_208_2; // @[Mux.scala 80:57]
  wire  _T_212_2 = _T_211 ? _T_2426 : _T_210_2; // @[Mux.scala 80:57]
  wire  _T_214_2 = _T_213 ? _T_2487 : _T_212_2; // @[Mux.scala 80:57]
  wire  _T_216_2 = _T_215 ? _T_2548 : _T_214_2; // @[Mux.scala 80:57]
  wire  _T_218_2 = _T_217 ? _T_2609 : _T_216_2; // @[Mux.scala 80:57]
  wire  _T_220_2 = _T_219 ? _T_2670 : _T_218_2; // @[Mux.scala 80:57]
  wire  _T_222_2 = _T_221 ? _T_2731 : _T_220_2; // @[Mux.scala 80:57]
  wire  _T_224_2 = _T_223 ? _T_2792 : _T_222_2; // @[Mux.scala 80:57]
  wire  _T_226_2 = _T_225 ? _T_2853 : _T_224_2; // @[Mux.scala 80:57]
  wire  _T_228_2 = _T_227 ? _T_2914 : _T_226_2; // @[Mux.scala 80:57]
  wire  _T_230_2 = _T_229 ? _T_2975 : _T_228_2; // @[Mux.scala 80:57]
  wire  _T_232_2 = _T_231 ? _T_3036 : _T_230_2; // @[Mux.scala 80:57]
  wire  _T_234_2 = _T_233 ? _T_3097 : _T_232_2; // @[Mux.scala 80:57]
  wire  _T_236_2 = _T_235 ? _T_3158 : _T_234_2; // @[Mux.scala 80:57]
  wire  _T_238_2 = _T_237 ? _T_3219 : _T_236_2; // @[Mux.scala 80:57]
  wire  _T_240_2 = _T_239 ? _T_3280 : _T_238_2; // @[Mux.scala 80:57]
  wire  _T_242_2 = _T_241 ? _T_3341 : _T_240_2; // @[Mux.scala 80:57]
  wire  _T_244_2 = _T_243 ? _T_3402 : _T_242_2; // @[Mux.scala 80:57]
  wire  _T_246_2 = _T_245 ? _T_3463 : _T_244_2; // @[Mux.scala 80:57]
  wire  _T_248_2 = _T_247 ? _T_3524 : _T_246_2; // @[Mux.scala 80:57]
  wire  _T_250_2 = _T_249 ? _T_3585 : _T_248_2; // @[Mux.scala 80:57]
  wire  _T_252_2 = _T_251 ? _T_3646 : _T_250_2; // @[Mux.scala 80:57]
  wire  _T_254_2 = _T_253 ? _T_3707 : _T_252_2; // @[Mux.scala 80:57]
  wire  _T_256_2 = _T_255 ? _T_3768 : _T_254_2; // @[Mux.scala 80:57]
  wire  _T_258_2 = _T_257 ? _T_3829 : _T_256_2; // @[Mux.scala 80:57]
  wire  _T_260_2 = _T_259 ? _T_3890 : _T_258_2; // @[Mux.scala 80:57]
  wire  _T_262_2 = _T_261 ? _T_3951 : _T_260_2; // @[Mux.scala 80:57]
  wire  _T_264_2 = _T_263 ? _T_4012 : _T_262_2; // @[Mux.scala 80:57]
  wire  _T_266_2 = _T_265 ? _T_4073 : _T_264_2; // @[Mux.scala 80:57]
  wire  _T_268_2 = _T_267 ? _T_4134 : _T_266_2; // @[Mux.scala 80:57]
  wire  _T_270_2 = _T_269 ? _T_4195 : _T_268_2; // @[Mux.scala 80:57]
  wire  _T_272_2 = _T_271 ? _T_4256 : _T_270_2; // @[Mux.scala 80:57]
  wire  _T_274_2 = _T_273 ? _T_4317 : _T_272_2; // @[Mux.scala 80:57]
  reg [21:0] _T_4309; // @[Reg.scala 27:20]
  reg [21:0] _T_4248; // @[Reg.scala 27:20]
  reg [21:0] _T_4187; // @[Reg.scala 27:20]
  reg [21:0] _T_4126; // @[Reg.scala 27:20]
  reg [21:0] _T_4065; // @[Reg.scala 27:20]
  reg [21:0] _T_4004; // @[Reg.scala 27:20]
  reg [21:0] _T_3943; // @[Reg.scala 27:20]
  reg [21:0] _T_3882; // @[Reg.scala 27:20]
  reg [21:0] _T_3821; // @[Reg.scala 27:20]
  reg [21:0] _T_3760; // @[Reg.scala 27:20]
  reg [21:0] _T_3699; // @[Reg.scala 27:20]
  reg [21:0] _T_3638; // @[Reg.scala 27:20]
  reg [21:0] _T_3577; // @[Reg.scala 27:20]
  reg [21:0] _T_3516; // @[Reg.scala 27:20]
  reg [21:0] _T_3455; // @[Reg.scala 27:20]
  reg [21:0] _T_3394; // @[Reg.scala 27:20]
  reg [21:0] _T_3333; // @[Reg.scala 27:20]
  reg [21:0] _T_3272; // @[Reg.scala 27:20]
  reg [21:0] _T_3211; // @[Reg.scala 27:20]
  reg [21:0] _T_3150; // @[Reg.scala 27:20]
  reg [21:0] _T_3089; // @[Reg.scala 27:20]
  reg [21:0] _T_3028; // @[Reg.scala 27:20]
  reg [21:0] _T_2967; // @[Reg.scala 27:20]
  reg [21:0] _T_2906; // @[Reg.scala 27:20]
  reg [21:0] _T_2845; // @[Reg.scala 27:20]
  reg [21:0] _T_2784; // @[Reg.scala 27:20]
  reg [21:0] _T_2723; // @[Reg.scala 27:20]
  reg [21:0] _T_2662; // @[Reg.scala 27:20]
  reg [21:0] _T_2601; // @[Reg.scala 27:20]
  reg [21:0] _T_2540; // @[Reg.scala 27:20]
  reg [21:0] _T_2479; // @[Reg.scala 27:20]
  reg [21:0] _T_2418; // @[Reg.scala 27:20]
  reg [21:0] _T_2357; // @[Reg.scala 27:20]
  reg [21:0] _T_2296; // @[Reg.scala 27:20]
  reg [21:0] _T_2235; // @[Reg.scala 27:20]
  reg [21:0] _T_2174; // @[Reg.scala 27:20]
  reg [21:0] _T_2113; // @[Reg.scala 27:20]
  reg [21:0] _T_2052; // @[Reg.scala 27:20]
  reg [21:0] _T_1991; // @[Reg.scala 27:20]
  reg [21:0] _T_1930; // @[Reg.scala 27:20]
  reg [21:0] _T_1869; // @[Reg.scala 27:20]
  reg [21:0] _T_1808; // @[Reg.scala 27:20]
  reg [21:0] _T_1747; // @[Reg.scala 27:20]
  reg [21:0] _T_1686; // @[Reg.scala 27:20]
  reg [21:0] _T_1625; // @[Reg.scala 27:20]
  reg [21:0] _T_1564; // @[Reg.scala 27:20]
  reg [21:0] _T_1503; // @[Reg.scala 27:20]
  reg [21:0] _T_1442; // @[Reg.scala 27:20]
  reg [21:0] _T_1381; // @[Reg.scala 27:20]
  reg [21:0] _T_1320; // @[Reg.scala 27:20]
  reg [21:0] _T_1259; // @[Reg.scala 27:20]
  reg [21:0] _T_1198; // @[Reg.scala 27:20]
  reg [21:0] _T_1137; // @[Reg.scala 27:20]
  reg [21:0] _T_1076; // @[Reg.scala 27:20]
  reg [21:0] _T_1015; // @[Reg.scala 27:20]
  reg [21:0] _T_954; // @[Reg.scala 27:20]
  reg [21:0] _T_893; // @[Reg.scala 27:20]
  reg [21:0] _T_832; // @[Reg.scala 27:20]
  reg [21:0] _T_771; // @[Reg.scala 27:20]
  reg [21:0] _T_710; // @[Reg.scala 27:20]
  reg [21:0] _T_649; // @[Reg.scala 27:20]
  reg [21:0] _T_588; // @[Reg.scala 27:20]
  reg [21:0] _T_527; // @[Reg.scala 27:20]
  reg [21:0] _T_466; // @[Reg.scala 27:20]
  wire [21:0] _T_24_2 = _T_149 ? _T_527 : _T_466; // @[Mux.scala 80:57]
  wire [21:0] _T_26_2 = _T_151 ? _T_588 : _T_24_2; // @[Mux.scala 80:57]
  wire [21:0] _T_28_2 = _T_153 ? _T_649 : _T_26_2; // @[Mux.scala 80:57]
  wire [21:0] _T_30_2 = _T_155 ? _T_710 : _T_28_2; // @[Mux.scala 80:57]
  wire [21:0] _T_32_2 = _T_157 ? _T_771 : _T_30_2; // @[Mux.scala 80:57]
  wire [21:0] _T_34_2 = _T_159 ? _T_832 : _T_32_2; // @[Mux.scala 80:57]
  wire [21:0] _T_36_2 = _T_161 ? _T_893 : _T_34_2; // @[Mux.scala 80:57]
  wire [21:0] _T_38_2 = _T_163 ? _T_954 : _T_36_2; // @[Mux.scala 80:57]
  wire [21:0] _T_40_2 = _T_165 ? _T_1015 : _T_38_2; // @[Mux.scala 80:57]
  wire [21:0] _T_42_2 = _T_167 ? _T_1076 : _T_40_2; // @[Mux.scala 80:57]
  wire [21:0] _T_44_2 = _T_169 ? _T_1137 : _T_42_2; // @[Mux.scala 80:57]
  wire [21:0] _T_46_2 = _T_171 ? _T_1198 : _T_44_2; // @[Mux.scala 80:57]
  wire [21:0] _T_48_2 = _T_173 ? _T_1259 : _T_46_2; // @[Mux.scala 80:57]
  wire [21:0] _T_50_2 = _T_175 ? _T_1320 : _T_48_2; // @[Mux.scala 80:57]
  wire [21:0] _T_52_2 = _T_177 ? _T_1381 : _T_50_2; // @[Mux.scala 80:57]
  wire [21:0] _T_54_2 = _T_179 ? _T_1442 : _T_52_2; // @[Mux.scala 80:57]
  wire [21:0] _T_56_2 = _T_181 ? _T_1503 : _T_54_2; // @[Mux.scala 80:57]
  wire [21:0] _T_58_2 = _T_183 ? _T_1564 : _T_56_2; // @[Mux.scala 80:57]
  wire [21:0] _T_60_2 = _T_185 ? _T_1625 : _T_58_2; // @[Mux.scala 80:57]
  wire [21:0] _T_62_2 = _T_187 ? _T_1686 : _T_60_2; // @[Mux.scala 80:57]
  wire [21:0] _T_64_2 = _T_189 ? _T_1747 : _T_62_2; // @[Mux.scala 80:57]
  wire [21:0] _T_66_2 = _T_191 ? _T_1808 : _T_64_2; // @[Mux.scala 80:57]
  wire [21:0] _T_68_2 = _T_193 ? _T_1869 : _T_66_2; // @[Mux.scala 80:57]
  wire [21:0] _T_70_2 = _T_195 ? _T_1930 : _T_68_2; // @[Mux.scala 80:57]
  wire [21:0] _T_72_2 = _T_197 ? _T_1991 : _T_70_2; // @[Mux.scala 80:57]
  wire [21:0] _T_74_2 = _T_199 ? _T_2052 : _T_72_2; // @[Mux.scala 80:57]
  wire [21:0] _T_76_2 = _T_201 ? _T_2113 : _T_74_2; // @[Mux.scala 80:57]
  wire [21:0] _T_78_2 = _T_203 ? _T_2174 : _T_76_2; // @[Mux.scala 80:57]
  wire [21:0] _T_80_2 = _T_205 ? _T_2235 : _T_78_2; // @[Mux.scala 80:57]
  wire [21:0] _T_82_2 = _T_207 ? _T_2296 : _T_80_2; // @[Mux.scala 80:57]
  wire [21:0] _T_84_2 = _T_209 ? _T_2357 : _T_82_2; // @[Mux.scala 80:57]
  wire [21:0] _T_86_2 = _T_211 ? _T_2418 : _T_84_2; // @[Mux.scala 80:57]
  wire [21:0] _T_88_2 = _T_213 ? _T_2479 : _T_86_2; // @[Mux.scala 80:57]
  wire [21:0] _T_90_2 = _T_215 ? _T_2540 : _T_88_2; // @[Mux.scala 80:57]
  wire [21:0] _T_92_2 = _T_217 ? _T_2601 : _T_90_2; // @[Mux.scala 80:57]
  wire [21:0] _T_94_2 = _T_219 ? _T_2662 : _T_92_2; // @[Mux.scala 80:57]
  wire [21:0] _T_96_2 = _T_221 ? _T_2723 : _T_94_2; // @[Mux.scala 80:57]
  wire [21:0] _T_98_2 = _T_223 ? _T_2784 : _T_96_2; // @[Mux.scala 80:57]
  wire [21:0] _T_100_2 = _T_225 ? _T_2845 : _T_98_2; // @[Mux.scala 80:57]
  wire [21:0] _T_102_2 = _T_227 ? _T_2906 : _T_100_2; // @[Mux.scala 80:57]
  wire [21:0] _T_104_2 = _T_229 ? _T_2967 : _T_102_2; // @[Mux.scala 80:57]
  wire [21:0] _T_106_2 = _T_231 ? _T_3028 : _T_104_2; // @[Mux.scala 80:57]
  wire [21:0] _T_108_2 = _T_233 ? _T_3089 : _T_106_2; // @[Mux.scala 80:57]
  wire [21:0] _T_110_2 = _T_235 ? _T_3150 : _T_108_2; // @[Mux.scala 80:57]
  wire [21:0] _T_112_2 = _T_237 ? _T_3211 : _T_110_2; // @[Mux.scala 80:57]
  wire [21:0] _T_114_2 = _T_239 ? _T_3272 : _T_112_2; // @[Mux.scala 80:57]
  wire [21:0] _T_116_2 = _T_241 ? _T_3333 : _T_114_2; // @[Mux.scala 80:57]
  wire [21:0] _T_118_2 = _T_243 ? _T_3394 : _T_116_2; // @[Mux.scala 80:57]
  wire [21:0] _T_120_2 = _T_245 ? _T_3455 : _T_118_2; // @[Mux.scala 80:57]
  wire [21:0] _T_122_2 = _T_247 ? _T_3516 : _T_120_2; // @[Mux.scala 80:57]
  wire [21:0] _T_124_2 = _T_249 ? _T_3577 : _T_122_2; // @[Mux.scala 80:57]
  wire [21:0] _T_126_2 = _T_251 ? _T_3638 : _T_124_2; // @[Mux.scala 80:57]
  wire [21:0] _T_128_2 = _T_253 ? _T_3699 : _T_126_2; // @[Mux.scala 80:57]
  wire [21:0] _T_130_2 = _T_255 ? _T_3760 : _T_128_2; // @[Mux.scala 80:57]
  wire [21:0] _T_132_2 = _T_257 ? _T_3821 : _T_130_2; // @[Mux.scala 80:57]
  wire [21:0] _T_134_2 = _T_259 ? _T_3882 : _T_132_2; // @[Mux.scala 80:57]
  wire [21:0] _T_136_2 = _T_261 ? _T_3943 : _T_134_2; // @[Mux.scala 80:57]
  wire [21:0] _T_138_2 = _T_263 ? _T_4004 : _T_136_2; // @[Mux.scala 80:57]
  wire [21:0] _T_140_2 = _T_265 ? _T_4065 : _T_138_2; // @[Mux.scala 80:57]
  wire [21:0] _T_142_2 = _T_267 ? _T_4126 : _T_140_2; // @[Mux.scala 80:57]
  wire [21:0] _T_144_2 = _T_269 ? _T_4187 : _T_142_2; // @[Mux.scala 80:57]
  wire [21:0] _T_146_2 = _T_271 ? _T_4248 : _T_144_2; // @[Mux.scala 80:57]
  wire [21:0] _T_148_2 = _T_273 ? _T_4309 : _T_146_2; // @[Mux.scala 80:57]
  wire  _T_279 = _T_148_2 == io_cacheIn_addr[31:10]; // @[Cache.scala 446:76]
  wire  _T_280 = _T_274_2 & _T_279; // @[Cache.scala 446:60]
  wire  _T_285 = _T_284 | _T_280; // @[Cache.scala 447:49]
  reg  _T_4331; // @[Reg.scala 27:20]
  reg  _T_4270; // @[Reg.scala 27:20]
  reg  _T_4209; // @[Reg.scala 27:20]
  reg  _T_4148; // @[Reg.scala 27:20]
  reg  _T_4087; // @[Reg.scala 27:20]
  reg  _T_4026; // @[Reg.scala 27:20]
  reg  _T_3965; // @[Reg.scala 27:20]
  reg  _T_3904; // @[Reg.scala 27:20]
  reg  _T_3843; // @[Reg.scala 27:20]
  reg  _T_3782; // @[Reg.scala 27:20]
  reg  _T_3721; // @[Reg.scala 27:20]
  reg  _T_3660; // @[Reg.scala 27:20]
  reg  _T_3599; // @[Reg.scala 27:20]
  reg  _T_3538; // @[Reg.scala 27:20]
  reg  _T_3477; // @[Reg.scala 27:20]
  reg  _T_3416; // @[Reg.scala 27:20]
  reg  _T_3355; // @[Reg.scala 27:20]
  reg  _T_3294; // @[Reg.scala 27:20]
  reg  _T_3233; // @[Reg.scala 27:20]
  reg  _T_3172; // @[Reg.scala 27:20]
  reg  _T_3111; // @[Reg.scala 27:20]
  reg  _T_3050; // @[Reg.scala 27:20]
  reg  _T_2989; // @[Reg.scala 27:20]
  reg  _T_2928; // @[Reg.scala 27:20]
  reg  _T_2867; // @[Reg.scala 27:20]
  reg  _T_2806; // @[Reg.scala 27:20]
  reg  _T_2745; // @[Reg.scala 27:20]
  reg  _T_2684; // @[Reg.scala 27:20]
  reg  _T_2623; // @[Reg.scala 27:20]
  reg  _T_2562; // @[Reg.scala 27:20]
  reg  _T_2501; // @[Reg.scala 27:20]
  reg  _T_2440; // @[Reg.scala 27:20]
  reg  _T_2379; // @[Reg.scala 27:20]
  reg  _T_2318; // @[Reg.scala 27:20]
  reg  _T_2257; // @[Reg.scala 27:20]
  reg  _T_2196; // @[Reg.scala 27:20]
  reg  _T_2135; // @[Reg.scala 27:20]
  reg  _T_2074; // @[Reg.scala 27:20]
  reg  _T_2013; // @[Reg.scala 27:20]
  reg  _T_1952; // @[Reg.scala 27:20]
  reg  _T_1891; // @[Reg.scala 27:20]
  reg  _T_1830; // @[Reg.scala 27:20]
  reg  _T_1769; // @[Reg.scala 27:20]
  reg  _T_1708; // @[Reg.scala 27:20]
  reg  _T_1647; // @[Reg.scala 27:20]
  reg  _T_1586; // @[Reg.scala 27:20]
  reg  _T_1525; // @[Reg.scala 27:20]
  reg  _T_1464; // @[Reg.scala 27:20]
  reg  _T_1403; // @[Reg.scala 27:20]
  reg  _T_1342; // @[Reg.scala 27:20]
  reg  _T_1281; // @[Reg.scala 27:20]
  reg  _T_1220; // @[Reg.scala 27:20]
  reg  _T_1159; // @[Reg.scala 27:20]
  reg  _T_1098; // @[Reg.scala 27:20]
  reg  _T_1037; // @[Reg.scala 27:20]
  reg  _T_976; // @[Reg.scala 27:20]
  reg  _T_915; // @[Reg.scala 27:20]
  reg  _T_854; // @[Reg.scala 27:20]
  reg  _T_793; // @[Reg.scala 27:20]
  reg  _T_732; // @[Reg.scala 27:20]
  reg  _T_671; // @[Reg.scala 27:20]
  reg  _T_610; // @[Reg.scala 27:20]
  reg  _T_549; // @[Reg.scala 27:20]
  reg  _T_488; // @[Reg.scala 27:20]
  wire  _T_150_3 = _T_149 ? _T_549 : _T_488; // @[Mux.scala 80:57]
  wire  _T_152_3 = _T_151 ? _T_610 : _T_150_3; // @[Mux.scala 80:57]
  wire  _T_154_3 = _T_153 ? _T_671 : _T_152_3; // @[Mux.scala 80:57]
  wire  _T_156_3 = _T_155 ? _T_732 : _T_154_3; // @[Mux.scala 80:57]
  wire  _T_158_3 = _T_157 ? _T_793 : _T_156_3; // @[Mux.scala 80:57]
  wire  _T_160_3 = _T_159 ? _T_854 : _T_158_3; // @[Mux.scala 80:57]
  wire  _T_162_3 = _T_161 ? _T_915 : _T_160_3; // @[Mux.scala 80:57]
  wire  _T_164_3 = _T_163 ? _T_976 : _T_162_3; // @[Mux.scala 80:57]
  wire  _T_166_3 = _T_165 ? _T_1037 : _T_164_3; // @[Mux.scala 80:57]
  wire  _T_168_3 = _T_167 ? _T_1098 : _T_166_3; // @[Mux.scala 80:57]
  wire  _T_170_3 = _T_169 ? _T_1159 : _T_168_3; // @[Mux.scala 80:57]
  wire  _T_172_3 = _T_171 ? _T_1220 : _T_170_3; // @[Mux.scala 80:57]
  wire  _T_174_3 = _T_173 ? _T_1281 : _T_172_3; // @[Mux.scala 80:57]
  wire  _T_176_3 = _T_175 ? _T_1342 : _T_174_3; // @[Mux.scala 80:57]
  wire  _T_178_3 = _T_177 ? _T_1403 : _T_176_3; // @[Mux.scala 80:57]
  wire  _T_180_3 = _T_179 ? _T_1464 : _T_178_3; // @[Mux.scala 80:57]
  wire  _T_182_3 = _T_181 ? _T_1525 : _T_180_3; // @[Mux.scala 80:57]
  wire  _T_184_3 = _T_183 ? _T_1586 : _T_182_3; // @[Mux.scala 80:57]
  wire  _T_186_3 = _T_185 ? _T_1647 : _T_184_3; // @[Mux.scala 80:57]
  wire  _T_188_3 = _T_187 ? _T_1708 : _T_186_3; // @[Mux.scala 80:57]
  wire  _T_190_3 = _T_189 ? _T_1769 : _T_188_3; // @[Mux.scala 80:57]
  wire  _T_192_3 = _T_191 ? _T_1830 : _T_190_3; // @[Mux.scala 80:57]
  wire  _T_194_3 = _T_193 ? _T_1891 : _T_192_3; // @[Mux.scala 80:57]
  wire  _T_196_3 = _T_195 ? _T_1952 : _T_194_3; // @[Mux.scala 80:57]
  wire  _T_198_3 = _T_197 ? _T_2013 : _T_196_3; // @[Mux.scala 80:57]
  wire  _T_200_3 = _T_199 ? _T_2074 : _T_198_3; // @[Mux.scala 80:57]
  wire  _T_202_3 = _T_201 ? _T_2135 : _T_200_3; // @[Mux.scala 80:57]
  wire  _T_204_3 = _T_203 ? _T_2196 : _T_202_3; // @[Mux.scala 80:57]
  wire  _T_206_3 = _T_205 ? _T_2257 : _T_204_3; // @[Mux.scala 80:57]
  wire  _T_208_3 = _T_207 ? _T_2318 : _T_206_3; // @[Mux.scala 80:57]
  wire  _T_210_3 = _T_209 ? _T_2379 : _T_208_3; // @[Mux.scala 80:57]
  wire  _T_212_3 = _T_211 ? _T_2440 : _T_210_3; // @[Mux.scala 80:57]
  wire  _T_214_3 = _T_213 ? _T_2501 : _T_212_3; // @[Mux.scala 80:57]
  wire  _T_216_3 = _T_215 ? _T_2562 : _T_214_3; // @[Mux.scala 80:57]
  wire  _T_218_3 = _T_217 ? _T_2623 : _T_216_3; // @[Mux.scala 80:57]
  wire  _T_220_3 = _T_219 ? _T_2684 : _T_218_3; // @[Mux.scala 80:57]
  wire  _T_222_3 = _T_221 ? _T_2745 : _T_220_3; // @[Mux.scala 80:57]
  wire  _T_224_3 = _T_223 ? _T_2806 : _T_222_3; // @[Mux.scala 80:57]
  wire  _T_226_3 = _T_225 ? _T_2867 : _T_224_3; // @[Mux.scala 80:57]
  wire  _T_228_3 = _T_227 ? _T_2928 : _T_226_3; // @[Mux.scala 80:57]
  wire  _T_230_3 = _T_229 ? _T_2989 : _T_228_3; // @[Mux.scala 80:57]
  wire  _T_232_3 = _T_231 ? _T_3050 : _T_230_3; // @[Mux.scala 80:57]
  wire  _T_234_3 = _T_233 ? _T_3111 : _T_232_3; // @[Mux.scala 80:57]
  wire  _T_236_3 = _T_235 ? _T_3172 : _T_234_3; // @[Mux.scala 80:57]
  wire  _T_238_3 = _T_237 ? _T_3233 : _T_236_3; // @[Mux.scala 80:57]
  wire  _T_240_3 = _T_239 ? _T_3294 : _T_238_3; // @[Mux.scala 80:57]
  wire  _T_242_3 = _T_241 ? _T_3355 : _T_240_3; // @[Mux.scala 80:57]
  wire  _T_244_3 = _T_243 ? _T_3416 : _T_242_3; // @[Mux.scala 80:57]
  wire  _T_246_3 = _T_245 ? _T_3477 : _T_244_3; // @[Mux.scala 80:57]
  wire  _T_248_3 = _T_247 ? _T_3538 : _T_246_3; // @[Mux.scala 80:57]
  wire  _T_250_3 = _T_249 ? _T_3599 : _T_248_3; // @[Mux.scala 80:57]
  wire  _T_252_3 = _T_251 ? _T_3660 : _T_250_3; // @[Mux.scala 80:57]
  wire  _T_254_3 = _T_253 ? _T_3721 : _T_252_3; // @[Mux.scala 80:57]
  wire  _T_256_3 = _T_255 ? _T_3782 : _T_254_3; // @[Mux.scala 80:57]
  wire  _T_258_3 = _T_257 ? _T_3843 : _T_256_3; // @[Mux.scala 80:57]
  wire  _T_260_3 = _T_259 ? _T_3904 : _T_258_3; // @[Mux.scala 80:57]
  wire  _T_262_3 = _T_261 ? _T_3965 : _T_260_3; // @[Mux.scala 80:57]
  wire  _T_264_3 = _T_263 ? _T_4026 : _T_262_3; // @[Mux.scala 80:57]
  wire  _T_266_3 = _T_265 ? _T_4087 : _T_264_3; // @[Mux.scala 80:57]
  wire  _T_268_3 = _T_267 ? _T_4148 : _T_266_3; // @[Mux.scala 80:57]
  wire  _T_270_3 = _T_269 ? _T_4209 : _T_268_3; // @[Mux.scala 80:57]
  wire  _T_272_3 = _T_271 ? _T_4270 : _T_270_3; // @[Mux.scala 80:57]
  wire  _T_274_3 = _T_273 ? _T_4331 : _T_272_3; // @[Mux.scala 80:57]
  reg [21:0] _T_4323; // @[Reg.scala 27:20]
  reg [21:0] _T_4262; // @[Reg.scala 27:20]
  reg [21:0] _T_4201; // @[Reg.scala 27:20]
  reg [21:0] _T_4140; // @[Reg.scala 27:20]
  reg [21:0] _T_4079; // @[Reg.scala 27:20]
  reg [21:0] _T_4018; // @[Reg.scala 27:20]
  reg [21:0] _T_3957; // @[Reg.scala 27:20]
  reg [21:0] _T_3896; // @[Reg.scala 27:20]
  reg [21:0] _T_3835; // @[Reg.scala 27:20]
  reg [21:0] _T_3774; // @[Reg.scala 27:20]
  reg [21:0] _T_3713; // @[Reg.scala 27:20]
  reg [21:0] _T_3652; // @[Reg.scala 27:20]
  reg [21:0] _T_3591; // @[Reg.scala 27:20]
  reg [21:0] _T_3530; // @[Reg.scala 27:20]
  reg [21:0] _T_3469; // @[Reg.scala 27:20]
  reg [21:0] _T_3408; // @[Reg.scala 27:20]
  reg [21:0] _T_3347; // @[Reg.scala 27:20]
  reg [21:0] _T_3286; // @[Reg.scala 27:20]
  reg [21:0] _T_3225; // @[Reg.scala 27:20]
  reg [21:0] _T_3164; // @[Reg.scala 27:20]
  reg [21:0] _T_3103; // @[Reg.scala 27:20]
  reg [21:0] _T_3042; // @[Reg.scala 27:20]
  reg [21:0] _T_2981; // @[Reg.scala 27:20]
  reg [21:0] _T_2920; // @[Reg.scala 27:20]
  reg [21:0] _T_2859; // @[Reg.scala 27:20]
  reg [21:0] _T_2798; // @[Reg.scala 27:20]
  reg [21:0] _T_2737; // @[Reg.scala 27:20]
  reg [21:0] _T_2676; // @[Reg.scala 27:20]
  reg [21:0] _T_2615; // @[Reg.scala 27:20]
  reg [21:0] _T_2554; // @[Reg.scala 27:20]
  reg [21:0] _T_2493; // @[Reg.scala 27:20]
  reg [21:0] _T_2432; // @[Reg.scala 27:20]
  reg [21:0] _T_2371; // @[Reg.scala 27:20]
  reg [21:0] _T_2310; // @[Reg.scala 27:20]
  reg [21:0] _T_2249; // @[Reg.scala 27:20]
  reg [21:0] _T_2188; // @[Reg.scala 27:20]
  reg [21:0] _T_2127; // @[Reg.scala 27:20]
  reg [21:0] _T_2066; // @[Reg.scala 27:20]
  reg [21:0] _T_2005; // @[Reg.scala 27:20]
  reg [21:0] _T_1944; // @[Reg.scala 27:20]
  reg [21:0] _T_1883; // @[Reg.scala 27:20]
  reg [21:0] _T_1822; // @[Reg.scala 27:20]
  reg [21:0] _T_1761; // @[Reg.scala 27:20]
  reg [21:0] _T_1700; // @[Reg.scala 27:20]
  reg [21:0] _T_1639; // @[Reg.scala 27:20]
  reg [21:0] _T_1578; // @[Reg.scala 27:20]
  reg [21:0] _T_1517; // @[Reg.scala 27:20]
  reg [21:0] _T_1456; // @[Reg.scala 27:20]
  reg [21:0] _T_1395; // @[Reg.scala 27:20]
  reg [21:0] _T_1334; // @[Reg.scala 27:20]
  reg [21:0] _T_1273; // @[Reg.scala 27:20]
  reg [21:0] _T_1212; // @[Reg.scala 27:20]
  reg [21:0] _T_1151; // @[Reg.scala 27:20]
  reg [21:0] _T_1090; // @[Reg.scala 27:20]
  reg [21:0] _T_1029; // @[Reg.scala 27:20]
  reg [21:0] _T_968; // @[Reg.scala 27:20]
  reg [21:0] _T_907; // @[Reg.scala 27:20]
  reg [21:0] _T_846; // @[Reg.scala 27:20]
  reg [21:0] _T_785; // @[Reg.scala 27:20]
  reg [21:0] _T_724; // @[Reg.scala 27:20]
  reg [21:0] _T_663; // @[Reg.scala 27:20]
  reg [21:0] _T_602; // @[Reg.scala 27:20]
  reg [21:0] _T_541; // @[Reg.scala 27:20]
  reg [21:0] _T_480; // @[Reg.scala 27:20]
  wire [21:0] _T_24_3 = _T_149 ? _T_541 : _T_480; // @[Mux.scala 80:57]
  wire [21:0] _T_26_3 = _T_151 ? _T_602 : _T_24_3; // @[Mux.scala 80:57]
  wire [21:0] _T_28_3 = _T_153 ? _T_663 : _T_26_3; // @[Mux.scala 80:57]
  wire [21:0] _T_30_3 = _T_155 ? _T_724 : _T_28_3; // @[Mux.scala 80:57]
  wire [21:0] _T_32_3 = _T_157 ? _T_785 : _T_30_3; // @[Mux.scala 80:57]
  wire [21:0] _T_34_3 = _T_159 ? _T_846 : _T_32_3; // @[Mux.scala 80:57]
  wire [21:0] _T_36_3 = _T_161 ? _T_907 : _T_34_3; // @[Mux.scala 80:57]
  wire [21:0] _T_38_3 = _T_163 ? _T_968 : _T_36_3; // @[Mux.scala 80:57]
  wire [21:0] _T_40_3 = _T_165 ? _T_1029 : _T_38_3; // @[Mux.scala 80:57]
  wire [21:0] _T_42_3 = _T_167 ? _T_1090 : _T_40_3; // @[Mux.scala 80:57]
  wire [21:0] _T_44_3 = _T_169 ? _T_1151 : _T_42_3; // @[Mux.scala 80:57]
  wire [21:0] _T_46_3 = _T_171 ? _T_1212 : _T_44_3; // @[Mux.scala 80:57]
  wire [21:0] _T_48_3 = _T_173 ? _T_1273 : _T_46_3; // @[Mux.scala 80:57]
  wire [21:0] _T_50_3 = _T_175 ? _T_1334 : _T_48_3; // @[Mux.scala 80:57]
  wire [21:0] _T_52_3 = _T_177 ? _T_1395 : _T_50_3; // @[Mux.scala 80:57]
  wire [21:0] _T_54_3 = _T_179 ? _T_1456 : _T_52_3; // @[Mux.scala 80:57]
  wire [21:0] _T_56_3 = _T_181 ? _T_1517 : _T_54_3; // @[Mux.scala 80:57]
  wire [21:0] _T_58_3 = _T_183 ? _T_1578 : _T_56_3; // @[Mux.scala 80:57]
  wire [21:0] _T_60_3 = _T_185 ? _T_1639 : _T_58_3; // @[Mux.scala 80:57]
  wire [21:0] _T_62_3 = _T_187 ? _T_1700 : _T_60_3; // @[Mux.scala 80:57]
  wire [21:0] _T_64_3 = _T_189 ? _T_1761 : _T_62_3; // @[Mux.scala 80:57]
  wire [21:0] _T_66_3 = _T_191 ? _T_1822 : _T_64_3; // @[Mux.scala 80:57]
  wire [21:0] _T_68_3 = _T_193 ? _T_1883 : _T_66_3; // @[Mux.scala 80:57]
  wire [21:0] _T_70_3 = _T_195 ? _T_1944 : _T_68_3; // @[Mux.scala 80:57]
  wire [21:0] _T_72_3 = _T_197 ? _T_2005 : _T_70_3; // @[Mux.scala 80:57]
  wire [21:0] _T_74_3 = _T_199 ? _T_2066 : _T_72_3; // @[Mux.scala 80:57]
  wire [21:0] _T_76_3 = _T_201 ? _T_2127 : _T_74_3; // @[Mux.scala 80:57]
  wire [21:0] _T_78_3 = _T_203 ? _T_2188 : _T_76_3; // @[Mux.scala 80:57]
  wire [21:0] _T_80_3 = _T_205 ? _T_2249 : _T_78_3; // @[Mux.scala 80:57]
  wire [21:0] _T_82_3 = _T_207 ? _T_2310 : _T_80_3; // @[Mux.scala 80:57]
  wire [21:0] _T_84_3 = _T_209 ? _T_2371 : _T_82_3; // @[Mux.scala 80:57]
  wire [21:0] _T_86_3 = _T_211 ? _T_2432 : _T_84_3; // @[Mux.scala 80:57]
  wire [21:0] _T_88_3 = _T_213 ? _T_2493 : _T_86_3; // @[Mux.scala 80:57]
  wire [21:0] _T_90_3 = _T_215 ? _T_2554 : _T_88_3; // @[Mux.scala 80:57]
  wire [21:0] _T_92_3 = _T_217 ? _T_2615 : _T_90_3; // @[Mux.scala 80:57]
  wire [21:0] _T_94_3 = _T_219 ? _T_2676 : _T_92_3; // @[Mux.scala 80:57]
  wire [21:0] _T_96_3 = _T_221 ? _T_2737 : _T_94_3; // @[Mux.scala 80:57]
  wire [21:0] _T_98_3 = _T_223 ? _T_2798 : _T_96_3; // @[Mux.scala 80:57]
  wire [21:0] _T_100_3 = _T_225 ? _T_2859 : _T_98_3; // @[Mux.scala 80:57]
  wire [21:0] _T_102_3 = _T_227 ? _T_2920 : _T_100_3; // @[Mux.scala 80:57]
  wire [21:0] _T_104_3 = _T_229 ? _T_2981 : _T_102_3; // @[Mux.scala 80:57]
  wire [21:0] _T_106_3 = _T_231 ? _T_3042 : _T_104_3; // @[Mux.scala 80:57]
  wire [21:0] _T_108_3 = _T_233 ? _T_3103 : _T_106_3; // @[Mux.scala 80:57]
  wire [21:0] _T_110_3 = _T_235 ? _T_3164 : _T_108_3; // @[Mux.scala 80:57]
  wire [21:0] _T_112_3 = _T_237 ? _T_3225 : _T_110_3; // @[Mux.scala 80:57]
  wire [21:0] _T_114_3 = _T_239 ? _T_3286 : _T_112_3; // @[Mux.scala 80:57]
  wire [21:0] _T_116_3 = _T_241 ? _T_3347 : _T_114_3; // @[Mux.scala 80:57]
  wire [21:0] _T_118_3 = _T_243 ? _T_3408 : _T_116_3; // @[Mux.scala 80:57]
  wire [21:0] _T_120_3 = _T_245 ? _T_3469 : _T_118_3; // @[Mux.scala 80:57]
  wire [21:0] _T_122_3 = _T_247 ? _T_3530 : _T_120_3; // @[Mux.scala 80:57]
  wire [21:0] _T_124_3 = _T_249 ? _T_3591 : _T_122_3; // @[Mux.scala 80:57]
  wire [21:0] _T_126_3 = _T_251 ? _T_3652 : _T_124_3; // @[Mux.scala 80:57]
  wire [21:0] _T_128_3 = _T_253 ? _T_3713 : _T_126_3; // @[Mux.scala 80:57]
  wire [21:0] _T_130_3 = _T_255 ? _T_3774 : _T_128_3; // @[Mux.scala 80:57]
  wire [21:0] _T_132_3 = _T_257 ? _T_3835 : _T_130_3; // @[Mux.scala 80:57]
  wire [21:0] _T_134_3 = _T_259 ? _T_3896 : _T_132_3; // @[Mux.scala 80:57]
  wire [21:0] _T_136_3 = _T_261 ? _T_3957 : _T_134_3; // @[Mux.scala 80:57]
  wire [21:0] _T_138_3 = _T_263 ? _T_4018 : _T_136_3; // @[Mux.scala 80:57]
  wire [21:0] _T_140_3 = _T_265 ? _T_4079 : _T_138_3; // @[Mux.scala 80:57]
  wire [21:0] _T_142_3 = _T_267 ? _T_4140 : _T_140_3; // @[Mux.scala 80:57]
  wire [21:0] _T_144_3 = _T_269 ? _T_4201 : _T_142_3; // @[Mux.scala 80:57]
  wire [21:0] _T_146_3 = _T_271 ? _T_4262 : _T_144_3; // @[Mux.scala 80:57]
  wire [21:0] _T_148_3 = _T_273 ? _T_4323 : _T_146_3; // @[Mux.scala 80:57]
  wire  _T_281 = _T_148_3 == io_cacheIn_addr[31:10]; // @[Cache.scala 446:76]
  wire  _T_282 = _T_274_3 & _T_281; // @[Cache.scala 446:60]
  wire  _T_286 = _T_285 | _T_282; // @[Cache.scala 447:49]
  wire  _T_11 = 2'h1 == _T_4; // @[Mux.scala 80:60]
  wire  _T_13 = 2'h2 == _T_4; // @[Mux.scala 80:60]
  wire  _T_15 = 2'h3 == _T_4; // @[Mux.scala 80:60]
  wire  _T_17 = _T_4 == 2'h0; // @[Cache.scala 417:27]
  wire  _T_18 = _T_4 == 2'h1; // @[Cache.scala 418:27]
  wire  _T_19 = _T_4 == 2'h2; // @[Cache.scala 419:27]
  wire  _T_20 = _T_4 == 2'h3; // @[Cache.scala 420:28]
  wire [127:0] _T_287 = _T_276 ? io_SRAMIO_0_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _T_288 = _T_278 ? io_SRAMIO_1_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _T_289 = _T_280 ? io_SRAMIO_2_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _T_290 = _T_282 ? io_SRAMIO_3_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _T_291 = _T_287 | _T_288; // @[Mux.scala 27:72]
  wire [127:0] _T_292 = _T_291 | _T_289; // @[Mux.scala 27:72]
  wire [127:0] _T_293 = _T_292 | _T_290; // @[Mux.scala 27:72]
  reg [1:0] _T_493; // @[Reg.scala 27:20]
  reg [1:0] _T_432; // @[Reg.scala 27:20]
  wire [1:0] _T_301 = _T_149 ? _T_493 : _T_432; // @[Mux.scala 80:57]
  reg [1:0] _T_554; // @[Reg.scala 27:20]
  wire [1:0] _T_303 = _T_151 ? _T_554 : _T_301; // @[Mux.scala 80:57]
  reg [1:0] _T_615; // @[Reg.scala 27:20]
  wire [1:0] _T_305 = _T_153 ? _T_615 : _T_303; // @[Mux.scala 80:57]
  reg [1:0] _T_676; // @[Reg.scala 27:20]
  wire [1:0] _T_307 = _T_155 ? _T_676 : _T_305; // @[Mux.scala 80:57]
  reg [1:0] _T_737; // @[Reg.scala 27:20]
  wire [1:0] _T_309 = _T_157 ? _T_737 : _T_307; // @[Mux.scala 80:57]
  reg [1:0] _T_798; // @[Reg.scala 27:20]
  wire [1:0] _T_311 = _T_159 ? _T_798 : _T_309; // @[Mux.scala 80:57]
  reg [1:0] _T_859; // @[Reg.scala 27:20]
  wire [1:0] _T_313 = _T_161 ? _T_859 : _T_311; // @[Mux.scala 80:57]
  reg [1:0] _T_920; // @[Reg.scala 27:20]
  wire [1:0] _T_315 = _T_163 ? _T_920 : _T_313; // @[Mux.scala 80:57]
  reg [1:0] _T_981; // @[Reg.scala 27:20]
  wire [1:0] _T_317 = _T_165 ? _T_981 : _T_315; // @[Mux.scala 80:57]
  reg [1:0] _T_1042; // @[Reg.scala 27:20]
  wire [1:0] _T_319 = _T_167 ? _T_1042 : _T_317; // @[Mux.scala 80:57]
  reg [1:0] _T_1103; // @[Reg.scala 27:20]
  wire [1:0] _T_321 = _T_169 ? _T_1103 : _T_319; // @[Mux.scala 80:57]
  reg [1:0] _T_1164; // @[Reg.scala 27:20]
  wire [1:0] _T_323 = _T_171 ? _T_1164 : _T_321; // @[Mux.scala 80:57]
  reg [1:0] _T_1225; // @[Reg.scala 27:20]
  wire [1:0] _T_325 = _T_173 ? _T_1225 : _T_323; // @[Mux.scala 80:57]
  reg [1:0] _T_1286; // @[Reg.scala 27:20]
  wire [1:0] _T_327 = _T_175 ? _T_1286 : _T_325; // @[Mux.scala 80:57]
  reg [1:0] _T_1347; // @[Reg.scala 27:20]
  wire [1:0] _T_329 = _T_177 ? _T_1347 : _T_327; // @[Mux.scala 80:57]
  reg [1:0] _T_1408; // @[Reg.scala 27:20]
  wire [1:0] _T_331 = _T_179 ? _T_1408 : _T_329; // @[Mux.scala 80:57]
  reg [1:0] _T_1469; // @[Reg.scala 27:20]
  wire [1:0] _T_333 = _T_181 ? _T_1469 : _T_331; // @[Mux.scala 80:57]
  reg [1:0] _T_1530; // @[Reg.scala 27:20]
  wire [1:0] _T_335 = _T_183 ? _T_1530 : _T_333; // @[Mux.scala 80:57]
  reg [1:0] _T_1591; // @[Reg.scala 27:20]
  wire [1:0] _T_337 = _T_185 ? _T_1591 : _T_335; // @[Mux.scala 80:57]
  reg [1:0] _T_1652; // @[Reg.scala 27:20]
  wire [1:0] _T_339 = _T_187 ? _T_1652 : _T_337; // @[Mux.scala 80:57]
  reg [1:0] _T_1713; // @[Reg.scala 27:20]
  wire [1:0] _T_341 = _T_189 ? _T_1713 : _T_339; // @[Mux.scala 80:57]
  reg [1:0] _T_1774; // @[Reg.scala 27:20]
  wire [1:0] _T_343 = _T_191 ? _T_1774 : _T_341; // @[Mux.scala 80:57]
  reg [1:0] _T_1835; // @[Reg.scala 27:20]
  wire [1:0] _T_345 = _T_193 ? _T_1835 : _T_343; // @[Mux.scala 80:57]
  reg [1:0] _T_1896; // @[Reg.scala 27:20]
  wire [1:0] _T_347 = _T_195 ? _T_1896 : _T_345; // @[Mux.scala 80:57]
  reg [1:0] _T_1957; // @[Reg.scala 27:20]
  wire [1:0] _T_349 = _T_197 ? _T_1957 : _T_347; // @[Mux.scala 80:57]
  reg [1:0] _T_2018; // @[Reg.scala 27:20]
  wire [1:0] _T_351 = _T_199 ? _T_2018 : _T_349; // @[Mux.scala 80:57]
  reg [1:0] _T_2079; // @[Reg.scala 27:20]
  wire [1:0] _T_353 = _T_201 ? _T_2079 : _T_351; // @[Mux.scala 80:57]
  reg [1:0] _T_2140; // @[Reg.scala 27:20]
  wire [1:0] _T_355 = _T_203 ? _T_2140 : _T_353; // @[Mux.scala 80:57]
  reg [1:0] _T_2201; // @[Reg.scala 27:20]
  wire [1:0] _T_357 = _T_205 ? _T_2201 : _T_355; // @[Mux.scala 80:57]
  reg [1:0] _T_2262; // @[Reg.scala 27:20]
  wire [1:0] _T_359 = _T_207 ? _T_2262 : _T_357; // @[Mux.scala 80:57]
  reg [1:0] _T_2323; // @[Reg.scala 27:20]
  wire [1:0] _T_361 = _T_209 ? _T_2323 : _T_359; // @[Mux.scala 80:57]
  reg [1:0] _T_2384; // @[Reg.scala 27:20]
  wire [1:0] _T_363 = _T_211 ? _T_2384 : _T_361; // @[Mux.scala 80:57]
  reg [1:0] _T_2445; // @[Reg.scala 27:20]
  wire [1:0] _T_365 = _T_213 ? _T_2445 : _T_363; // @[Mux.scala 80:57]
  reg [1:0] _T_2506; // @[Reg.scala 27:20]
  wire [1:0] _T_367 = _T_215 ? _T_2506 : _T_365; // @[Mux.scala 80:57]
  reg [1:0] _T_2567; // @[Reg.scala 27:20]
  wire [1:0] _T_369 = _T_217 ? _T_2567 : _T_367; // @[Mux.scala 80:57]
  reg [1:0] _T_2628; // @[Reg.scala 27:20]
  wire [1:0] _T_371 = _T_219 ? _T_2628 : _T_369; // @[Mux.scala 80:57]
  reg [1:0] _T_2689; // @[Reg.scala 27:20]
  wire [1:0] _T_373 = _T_221 ? _T_2689 : _T_371; // @[Mux.scala 80:57]
  reg [1:0] _T_2750; // @[Reg.scala 27:20]
  wire [1:0] _T_375 = _T_223 ? _T_2750 : _T_373; // @[Mux.scala 80:57]
  reg [1:0] _T_2811; // @[Reg.scala 27:20]
  wire [1:0] _T_377 = _T_225 ? _T_2811 : _T_375; // @[Mux.scala 80:57]
  reg [1:0] _T_2872; // @[Reg.scala 27:20]
  wire [1:0] _T_379 = _T_227 ? _T_2872 : _T_377; // @[Mux.scala 80:57]
  reg [1:0] _T_2933; // @[Reg.scala 27:20]
  wire [1:0] _T_381 = _T_229 ? _T_2933 : _T_379; // @[Mux.scala 80:57]
  reg [1:0] _T_2994; // @[Reg.scala 27:20]
  wire [1:0] _T_383 = _T_231 ? _T_2994 : _T_381; // @[Mux.scala 80:57]
  reg [1:0] _T_3055; // @[Reg.scala 27:20]
  wire [1:0] _T_385 = _T_233 ? _T_3055 : _T_383; // @[Mux.scala 80:57]
  reg [1:0] _T_3116; // @[Reg.scala 27:20]
  wire [1:0] _T_387 = _T_235 ? _T_3116 : _T_385; // @[Mux.scala 80:57]
  reg [1:0] _T_3177; // @[Reg.scala 27:20]
  wire [1:0] _T_389 = _T_237 ? _T_3177 : _T_387; // @[Mux.scala 80:57]
  reg [1:0] _T_3238; // @[Reg.scala 27:20]
  wire [1:0] _T_391 = _T_239 ? _T_3238 : _T_389; // @[Mux.scala 80:57]
  reg [1:0] _T_3299; // @[Reg.scala 27:20]
  wire [1:0] _T_393 = _T_241 ? _T_3299 : _T_391; // @[Mux.scala 80:57]
  reg [1:0] _T_3360; // @[Reg.scala 27:20]
  wire [1:0] _T_395 = _T_243 ? _T_3360 : _T_393; // @[Mux.scala 80:57]
  reg [1:0] _T_3421; // @[Reg.scala 27:20]
  wire [1:0] _T_397 = _T_245 ? _T_3421 : _T_395; // @[Mux.scala 80:57]
  reg [1:0] _T_3482; // @[Reg.scala 27:20]
  wire [1:0] _T_399 = _T_247 ? _T_3482 : _T_397; // @[Mux.scala 80:57]
  reg [1:0] _T_3543; // @[Reg.scala 27:20]
  wire [1:0] _T_401 = _T_249 ? _T_3543 : _T_399; // @[Mux.scala 80:57]
  reg [1:0] _T_3604; // @[Reg.scala 27:20]
  wire [1:0] _T_403 = _T_251 ? _T_3604 : _T_401; // @[Mux.scala 80:57]
  reg [1:0] _T_3665; // @[Reg.scala 27:20]
  wire [1:0] _T_405 = _T_253 ? _T_3665 : _T_403; // @[Mux.scala 80:57]
  reg [1:0] _T_3726; // @[Reg.scala 27:20]
  wire [1:0] _T_407 = _T_255 ? _T_3726 : _T_405; // @[Mux.scala 80:57]
  reg [1:0] _T_3787; // @[Reg.scala 27:20]
  wire [1:0] _T_409 = _T_257 ? _T_3787 : _T_407; // @[Mux.scala 80:57]
  reg [1:0] _T_3848; // @[Reg.scala 27:20]
  wire [1:0] _T_411 = _T_259 ? _T_3848 : _T_409; // @[Mux.scala 80:57]
  reg [1:0] _T_3909; // @[Reg.scala 27:20]
  wire [1:0] _T_413 = _T_261 ? _T_3909 : _T_411; // @[Mux.scala 80:57]
  reg [1:0] _T_3970; // @[Reg.scala 27:20]
  wire [1:0] _T_415 = _T_263 ? _T_3970 : _T_413; // @[Mux.scala 80:57]
  reg [1:0] _T_4031; // @[Reg.scala 27:20]
  wire [1:0] _T_417 = _T_265 ? _T_4031 : _T_415; // @[Mux.scala 80:57]
  reg [1:0] _T_4092; // @[Reg.scala 27:20]
  wire [1:0] _T_419 = _T_267 ? _T_4092 : _T_417; // @[Mux.scala 80:57]
  reg [1:0] _T_4153; // @[Reg.scala 27:20]
  wire [1:0] _T_421 = _T_269 ? _T_4153 : _T_419; // @[Mux.scala 80:57]
  reg [1:0] _T_4214; // @[Reg.scala 27:20]
  wire [1:0] _T_423 = _T_271 ? _T_4214 : _T_421; // @[Mux.scala 80:57]
  reg [1:0] _T_4275; // @[Reg.scala 27:20]
  wire [1:0] _T_425 = _T_273 ? _T_4275 : _T_423; // @[Mux.scala 80:57]
  wire [1:0] _T_429 = _T_432 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_430 = 6'h0 == io_cacheIn_addr[9:4]; // @[Cache.scala 488:35]
  wire  _T_431 = io_cacheOut_r_last_i & _T_430; // @[Cache.scala 488:28]
  wire  _T_435 = _T_432 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_436 = _T_431 & _T_435; // @[Cache.scala 491:87]
  wire  _T_437 = _T_436 & _T_18; // @[Cache.scala 491:114]
  wire  _T_440 = reset | updataICache; // @[Cache.scala 492:32]
  wire  _GEN_2 = _T_437 | _T_446; // @[Reg.scala 28:19]
  wire  _T_449 = _T_432 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_450 = _T_431 & _T_449; // @[Cache.scala 491:87]
  wire  _T_451 = _T_450 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_4 = _T_451 | _T_460; // @[Reg.scala 28:19]
  wire  _T_463 = _T_432 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_464 = _T_431 & _T_463; // @[Cache.scala 491:87]
  wire  _T_465 = _T_464 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_6 = _T_465 | _T_474; // @[Reg.scala 28:19]
  wire  _T_477 = _T_432 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_478 = _T_431 & _T_477; // @[Cache.scala 491:87]
  wire  _T_479 = _T_478 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_8 = _T_479 | _T_488; // @[Reg.scala 28:19]
  wire [1:0] _T_490 = _T_493 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_492 = io_cacheOut_r_last_i & _T_149; // @[Cache.scala 488:28]
  wire  _T_496 = _T_493 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_497 = _T_492 & _T_496; // @[Cache.scala 491:87]
  wire  _T_498 = _T_497 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_11 = _T_498 | _T_507; // @[Reg.scala 28:19]
  wire  _T_510 = _T_493 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_511 = _T_492 & _T_510; // @[Cache.scala 491:87]
  wire  _T_512 = _T_511 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_13 = _T_512 | _T_521; // @[Reg.scala 28:19]
  wire  _T_524 = _T_493 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_525 = _T_492 & _T_524; // @[Cache.scala 491:87]
  wire  _T_526 = _T_525 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_15 = _T_526 | _T_535; // @[Reg.scala 28:19]
  wire  _T_538 = _T_493 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_539 = _T_492 & _T_538; // @[Cache.scala 491:87]
  wire  _T_540 = _T_539 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_17 = _T_540 | _T_549; // @[Reg.scala 28:19]
  wire [1:0] _T_551 = _T_554 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_553 = io_cacheOut_r_last_i & _T_151; // @[Cache.scala 488:28]
  wire  _T_557 = _T_554 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_558 = _T_553 & _T_557; // @[Cache.scala 491:87]
  wire  _T_559 = _T_558 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_20 = _T_559 | _T_568; // @[Reg.scala 28:19]
  wire  _T_571 = _T_554 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_572 = _T_553 & _T_571; // @[Cache.scala 491:87]
  wire  _T_573 = _T_572 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_22 = _T_573 | _T_582; // @[Reg.scala 28:19]
  wire  _T_585 = _T_554 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_586 = _T_553 & _T_585; // @[Cache.scala 491:87]
  wire  _T_587 = _T_586 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_24 = _T_587 | _T_596; // @[Reg.scala 28:19]
  wire  _T_599 = _T_554 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_600 = _T_553 & _T_599; // @[Cache.scala 491:87]
  wire  _T_601 = _T_600 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_26 = _T_601 | _T_610; // @[Reg.scala 28:19]
  wire [1:0] _T_612 = _T_615 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_614 = io_cacheOut_r_last_i & _T_153; // @[Cache.scala 488:28]
  wire  _T_618 = _T_615 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_619 = _T_614 & _T_618; // @[Cache.scala 491:87]
  wire  _T_620 = _T_619 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_29 = _T_620 | _T_629; // @[Reg.scala 28:19]
  wire  _T_632 = _T_615 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_633 = _T_614 & _T_632; // @[Cache.scala 491:87]
  wire  _T_634 = _T_633 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_31 = _T_634 | _T_643; // @[Reg.scala 28:19]
  wire  _T_646 = _T_615 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_647 = _T_614 & _T_646; // @[Cache.scala 491:87]
  wire  _T_648 = _T_647 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_33 = _T_648 | _T_657; // @[Reg.scala 28:19]
  wire  _T_660 = _T_615 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_661 = _T_614 & _T_660; // @[Cache.scala 491:87]
  wire  _T_662 = _T_661 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_35 = _T_662 | _T_671; // @[Reg.scala 28:19]
  wire [1:0] _T_673 = _T_676 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_675 = io_cacheOut_r_last_i & _T_155; // @[Cache.scala 488:28]
  wire  _T_679 = _T_676 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_680 = _T_675 & _T_679; // @[Cache.scala 491:87]
  wire  _T_681 = _T_680 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_38 = _T_681 | _T_690; // @[Reg.scala 28:19]
  wire  _T_693 = _T_676 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_694 = _T_675 & _T_693; // @[Cache.scala 491:87]
  wire  _T_695 = _T_694 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_40 = _T_695 | _T_704; // @[Reg.scala 28:19]
  wire  _T_707 = _T_676 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_708 = _T_675 & _T_707; // @[Cache.scala 491:87]
  wire  _T_709 = _T_708 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_42 = _T_709 | _T_718; // @[Reg.scala 28:19]
  wire  _T_721 = _T_676 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_722 = _T_675 & _T_721; // @[Cache.scala 491:87]
  wire  _T_723 = _T_722 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_44 = _T_723 | _T_732; // @[Reg.scala 28:19]
  wire [1:0] _T_734 = _T_737 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_736 = io_cacheOut_r_last_i & _T_157; // @[Cache.scala 488:28]
  wire  _T_740 = _T_737 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_741 = _T_736 & _T_740; // @[Cache.scala 491:87]
  wire  _T_742 = _T_741 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_47 = _T_742 | _T_751; // @[Reg.scala 28:19]
  wire  _T_754 = _T_737 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_755 = _T_736 & _T_754; // @[Cache.scala 491:87]
  wire  _T_756 = _T_755 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_49 = _T_756 | _T_765; // @[Reg.scala 28:19]
  wire  _T_768 = _T_737 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_769 = _T_736 & _T_768; // @[Cache.scala 491:87]
  wire  _T_770 = _T_769 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_51 = _T_770 | _T_779; // @[Reg.scala 28:19]
  wire  _T_782 = _T_737 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_783 = _T_736 & _T_782; // @[Cache.scala 491:87]
  wire  _T_784 = _T_783 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_53 = _T_784 | _T_793; // @[Reg.scala 28:19]
  wire [1:0] _T_795 = _T_798 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_797 = io_cacheOut_r_last_i & _T_159; // @[Cache.scala 488:28]
  wire  _T_801 = _T_798 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_802 = _T_797 & _T_801; // @[Cache.scala 491:87]
  wire  _T_803 = _T_802 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_56 = _T_803 | _T_812; // @[Reg.scala 28:19]
  wire  _T_815 = _T_798 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_816 = _T_797 & _T_815; // @[Cache.scala 491:87]
  wire  _T_817 = _T_816 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_58 = _T_817 | _T_826; // @[Reg.scala 28:19]
  wire  _T_829 = _T_798 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_830 = _T_797 & _T_829; // @[Cache.scala 491:87]
  wire  _T_831 = _T_830 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_60 = _T_831 | _T_840; // @[Reg.scala 28:19]
  wire  _T_843 = _T_798 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_844 = _T_797 & _T_843; // @[Cache.scala 491:87]
  wire  _T_845 = _T_844 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_62 = _T_845 | _T_854; // @[Reg.scala 28:19]
  wire [1:0] _T_856 = _T_859 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_858 = io_cacheOut_r_last_i & _T_161; // @[Cache.scala 488:28]
  wire  _T_862 = _T_859 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_863 = _T_858 & _T_862; // @[Cache.scala 491:87]
  wire  _T_864 = _T_863 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_65 = _T_864 | _T_873; // @[Reg.scala 28:19]
  wire  _T_876 = _T_859 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_877 = _T_858 & _T_876; // @[Cache.scala 491:87]
  wire  _T_878 = _T_877 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_67 = _T_878 | _T_887; // @[Reg.scala 28:19]
  wire  _T_890 = _T_859 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_891 = _T_858 & _T_890; // @[Cache.scala 491:87]
  wire  _T_892 = _T_891 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_69 = _T_892 | _T_901; // @[Reg.scala 28:19]
  wire  _T_904 = _T_859 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_905 = _T_858 & _T_904; // @[Cache.scala 491:87]
  wire  _T_906 = _T_905 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_71 = _T_906 | _T_915; // @[Reg.scala 28:19]
  wire [1:0] _T_917 = _T_920 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_919 = io_cacheOut_r_last_i & _T_163; // @[Cache.scala 488:28]
  wire  _T_923 = _T_920 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_924 = _T_919 & _T_923; // @[Cache.scala 491:87]
  wire  _T_925 = _T_924 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_74 = _T_925 | _T_934; // @[Reg.scala 28:19]
  wire  _T_937 = _T_920 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_938 = _T_919 & _T_937; // @[Cache.scala 491:87]
  wire  _T_939 = _T_938 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_76 = _T_939 | _T_948; // @[Reg.scala 28:19]
  wire  _T_951 = _T_920 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_952 = _T_919 & _T_951; // @[Cache.scala 491:87]
  wire  _T_953 = _T_952 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_78 = _T_953 | _T_962; // @[Reg.scala 28:19]
  wire  _T_965 = _T_920 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_966 = _T_919 & _T_965; // @[Cache.scala 491:87]
  wire  _T_967 = _T_966 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_80 = _T_967 | _T_976; // @[Reg.scala 28:19]
  wire [1:0] _T_978 = _T_981 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_980 = io_cacheOut_r_last_i & _T_165; // @[Cache.scala 488:28]
  wire  _T_984 = _T_981 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_985 = _T_980 & _T_984; // @[Cache.scala 491:87]
  wire  _T_986 = _T_985 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_83 = _T_986 | _T_995; // @[Reg.scala 28:19]
  wire  _T_998 = _T_981 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_999 = _T_980 & _T_998; // @[Cache.scala 491:87]
  wire  _T_1000 = _T_999 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_85 = _T_1000 | _T_1009; // @[Reg.scala 28:19]
  wire  _T_1012 = _T_981 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_1013 = _T_980 & _T_1012; // @[Cache.scala 491:87]
  wire  _T_1014 = _T_1013 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_87 = _T_1014 | _T_1023; // @[Reg.scala 28:19]
  wire  _T_1026 = _T_981 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_1027 = _T_980 & _T_1026; // @[Cache.scala 491:87]
  wire  _T_1028 = _T_1027 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_89 = _T_1028 | _T_1037; // @[Reg.scala 28:19]
  wire [1:0] _T_1039 = _T_1042 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_1041 = io_cacheOut_r_last_i & _T_167; // @[Cache.scala 488:28]
  wire  _T_1045 = _T_1042 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_1046 = _T_1041 & _T_1045; // @[Cache.scala 491:87]
  wire  _T_1047 = _T_1046 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_92 = _T_1047 | _T_1056; // @[Reg.scala 28:19]
  wire  _T_1059 = _T_1042 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_1060 = _T_1041 & _T_1059; // @[Cache.scala 491:87]
  wire  _T_1061 = _T_1060 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_94 = _T_1061 | _T_1070; // @[Reg.scala 28:19]
  wire  _T_1073 = _T_1042 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_1074 = _T_1041 & _T_1073; // @[Cache.scala 491:87]
  wire  _T_1075 = _T_1074 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_96 = _T_1075 | _T_1084; // @[Reg.scala 28:19]
  wire  _T_1087 = _T_1042 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_1088 = _T_1041 & _T_1087; // @[Cache.scala 491:87]
  wire  _T_1089 = _T_1088 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_98 = _T_1089 | _T_1098; // @[Reg.scala 28:19]
  wire [1:0] _T_1100 = _T_1103 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_1102 = io_cacheOut_r_last_i & _T_169; // @[Cache.scala 488:28]
  wire  _T_1106 = _T_1103 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_1107 = _T_1102 & _T_1106; // @[Cache.scala 491:87]
  wire  _T_1108 = _T_1107 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_101 = _T_1108 | _T_1117; // @[Reg.scala 28:19]
  wire  _T_1120 = _T_1103 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_1121 = _T_1102 & _T_1120; // @[Cache.scala 491:87]
  wire  _T_1122 = _T_1121 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_103 = _T_1122 | _T_1131; // @[Reg.scala 28:19]
  wire  _T_1134 = _T_1103 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_1135 = _T_1102 & _T_1134; // @[Cache.scala 491:87]
  wire  _T_1136 = _T_1135 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_105 = _T_1136 | _T_1145; // @[Reg.scala 28:19]
  wire  _T_1148 = _T_1103 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_1149 = _T_1102 & _T_1148; // @[Cache.scala 491:87]
  wire  _T_1150 = _T_1149 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_107 = _T_1150 | _T_1159; // @[Reg.scala 28:19]
  wire [1:0] _T_1161 = _T_1164 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_1163 = io_cacheOut_r_last_i & _T_171; // @[Cache.scala 488:28]
  wire  _T_1167 = _T_1164 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_1168 = _T_1163 & _T_1167; // @[Cache.scala 491:87]
  wire  _T_1169 = _T_1168 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_110 = _T_1169 | _T_1178; // @[Reg.scala 28:19]
  wire  _T_1181 = _T_1164 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_1182 = _T_1163 & _T_1181; // @[Cache.scala 491:87]
  wire  _T_1183 = _T_1182 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_112 = _T_1183 | _T_1192; // @[Reg.scala 28:19]
  wire  _T_1195 = _T_1164 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_1196 = _T_1163 & _T_1195; // @[Cache.scala 491:87]
  wire  _T_1197 = _T_1196 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_114 = _T_1197 | _T_1206; // @[Reg.scala 28:19]
  wire  _T_1209 = _T_1164 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_1210 = _T_1163 & _T_1209; // @[Cache.scala 491:87]
  wire  _T_1211 = _T_1210 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_116 = _T_1211 | _T_1220; // @[Reg.scala 28:19]
  wire [1:0] _T_1222 = _T_1225 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_1224 = io_cacheOut_r_last_i & _T_173; // @[Cache.scala 488:28]
  wire  _T_1228 = _T_1225 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_1229 = _T_1224 & _T_1228; // @[Cache.scala 491:87]
  wire  _T_1230 = _T_1229 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_119 = _T_1230 | _T_1239; // @[Reg.scala 28:19]
  wire  _T_1242 = _T_1225 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_1243 = _T_1224 & _T_1242; // @[Cache.scala 491:87]
  wire  _T_1244 = _T_1243 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_121 = _T_1244 | _T_1253; // @[Reg.scala 28:19]
  wire  _T_1256 = _T_1225 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_1257 = _T_1224 & _T_1256; // @[Cache.scala 491:87]
  wire  _T_1258 = _T_1257 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_123 = _T_1258 | _T_1267; // @[Reg.scala 28:19]
  wire  _T_1270 = _T_1225 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_1271 = _T_1224 & _T_1270; // @[Cache.scala 491:87]
  wire  _T_1272 = _T_1271 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_125 = _T_1272 | _T_1281; // @[Reg.scala 28:19]
  wire [1:0] _T_1283 = _T_1286 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_1285 = io_cacheOut_r_last_i & _T_175; // @[Cache.scala 488:28]
  wire  _T_1289 = _T_1286 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_1290 = _T_1285 & _T_1289; // @[Cache.scala 491:87]
  wire  _T_1291 = _T_1290 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_128 = _T_1291 | _T_1300; // @[Reg.scala 28:19]
  wire  _T_1303 = _T_1286 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_1304 = _T_1285 & _T_1303; // @[Cache.scala 491:87]
  wire  _T_1305 = _T_1304 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_130 = _T_1305 | _T_1314; // @[Reg.scala 28:19]
  wire  _T_1317 = _T_1286 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_1318 = _T_1285 & _T_1317; // @[Cache.scala 491:87]
  wire  _T_1319 = _T_1318 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_132 = _T_1319 | _T_1328; // @[Reg.scala 28:19]
  wire  _T_1331 = _T_1286 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_1332 = _T_1285 & _T_1331; // @[Cache.scala 491:87]
  wire  _T_1333 = _T_1332 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_134 = _T_1333 | _T_1342; // @[Reg.scala 28:19]
  wire [1:0] _T_1344 = _T_1347 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_1346 = io_cacheOut_r_last_i & _T_177; // @[Cache.scala 488:28]
  wire  _T_1350 = _T_1347 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_1351 = _T_1346 & _T_1350; // @[Cache.scala 491:87]
  wire  _T_1352 = _T_1351 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_137 = _T_1352 | _T_1361; // @[Reg.scala 28:19]
  wire  _T_1364 = _T_1347 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_1365 = _T_1346 & _T_1364; // @[Cache.scala 491:87]
  wire  _T_1366 = _T_1365 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_139 = _T_1366 | _T_1375; // @[Reg.scala 28:19]
  wire  _T_1378 = _T_1347 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_1379 = _T_1346 & _T_1378; // @[Cache.scala 491:87]
  wire  _T_1380 = _T_1379 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_141 = _T_1380 | _T_1389; // @[Reg.scala 28:19]
  wire  _T_1392 = _T_1347 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_1393 = _T_1346 & _T_1392; // @[Cache.scala 491:87]
  wire  _T_1394 = _T_1393 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_143 = _T_1394 | _T_1403; // @[Reg.scala 28:19]
  wire [1:0] _T_1405 = _T_1408 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_1407 = io_cacheOut_r_last_i & _T_179; // @[Cache.scala 488:28]
  wire  _T_1411 = _T_1408 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_1412 = _T_1407 & _T_1411; // @[Cache.scala 491:87]
  wire  _T_1413 = _T_1412 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_146 = _T_1413 | _T_1422; // @[Reg.scala 28:19]
  wire  _T_1425 = _T_1408 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_1426 = _T_1407 & _T_1425; // @[Cache.scala 491:87]
  wire  _T_1427 = _T_1426 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_148 = _T_1427 | _T_1436; // @[Reg.scala 28:19]
  wire  _T_1439 = _T_1408 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_1440 = _T_1407 & _T_1439; // @[Cache.scala 491:87]
  wire  _T_1441 = _T_1440 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_150 = _T_1441 | _T_1450; // @[Reg.scala 28:19]
  wire  _T_1453 = _T_1408 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_1454 = _T_1407 & _T_1453; // @[Cache.scala 491:87]
  wire  _T_1455 = _T_1454 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_152 = _T_1455 | _T_1464; // @[Reg.scala 28:19]
  wire [1:0] _T_1466 = _T_1469 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_1468 = io_cacheOut_r_last_i & _T_181; // @[Cache.scala 488:28]
  wire  _T_1472 = _T_1469 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_1473 = _T_1468 & _T_1472; // @[Cache.scala 491:87]
  wire  _T_1474 = _T_1473 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_155 = _T_1474 | _T_1483; // @[Reg.scala 28:19]
  wire  _T_1486 = _T_1469 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_1487 = _T_1468 & _T_1486; // @[Cache.scala 491:87]
  wire  _T_1488 = _T_1487 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_157 = _T_1488 | _T_1497; // @[Reg.scala 28:19]
  wire  _T_1500 = _T_1469 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_1501 = _T_1468 & _T_1500; // @[Cache.scala 491:87]
  wire  _T_1502 = _T_1501 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_159 = _T_1502 | _T_1511; // @[Reg.scala 28:19]
  wire  _T_1514 = _T_1469 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_1515 = _T_1468 & _T_1514; // @[Cache.scala 491:87]
  wire  _T_1516 = _T_1515 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_161 = _T_1516 | _T_1525; // @[Reg.scala 28:19]
  wire [1:0] _T_1527 = _T_1530 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_1529 = io_cacheOut_r_last_i & _T_183; // @[Cache.scala 488:28]
  wire  _T_1533 = _T_1530 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_1534 = _T_1529 & _T_1533; // @[Cache.scala 491:87]
  wire  _T_1535 = _T_1534 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_164 = _T_1535 | _T_1544; // @[Reg.scala 28:19]
  wire  _T_1547 = _T_1530 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_1548 = _T_1529 & _T_1547; // @[Cache.scala 491:87]
  wire  _T_1549 = _T_1548 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_166 = _T_1549 | _T_1558; // @[Reg.scala 28:19]
  wire  _T_1561 = _T_1530 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_1562 = _T_1529 & _T_1561; // @[Cache.scala 491:87]
  wire  _T_1563 = _T_1562 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_168 = _T_1563 | _T_1572; // @[Reg.scala 28:19]
  wire  _T_1575 = _T_1530 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_1576 = _T_1529 & _T_1575; // @[Cache.scala 491:87]
  wire  _T_1577 = _T_1576 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_170 = _T_1577 | _T_1586; // @[Reg.scala 28:19]
  wire [1:0] _T_1588 = _T_1591 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_1590 = io_cacheOut_r_last_i & _T_185; // @[Cache.scala 488:28]
  wire  _T_1594 = _T_1591 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_1595 = _T_1590 & _T_1594; // @[Cache.scala 491:87]
  wire  _T_1596 = _T_1595 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_173 = _T_1596 | _T_1605; // @[Reg.scala 28:19]
  wire  _T_1608 = _T_1591 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_1609 = _T_1590 & _T_1608; // @[Cache.scala 491:87]
  wire  _T_1610 = _T_1609 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_175 = _T_1610 | _T_1619; // @[Reg.scala 28:19]
  wire  _T_1622 = _T_1591 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_1623 = _T_1590 & _T_1622; // @[Cache.scala 491:87]
  wire  _T_1624 = _T_1623 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_177 = _T_1624 | _T_1633; // @[Reg.scala 28:19]
  wire  _T_1636 = _T_1591 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_1637 = _T_1590 & _T_1636; // @[Cache.scala 491:87]
  wire  _T_1638 = _T_1637 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_179 = _T_1638 | _T_1647; // @[Reg.scala 28:19]
  wire [1:0] _T_1649 = _T_1652 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_1651 = io_cacheOut_r_last_i & _T_187; // @[Cache.scala 488:28]
  wire  _T_1655 = _T_1652 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_1656 = _T_1651 & _T_1655; // @[Cache.scala 491:87]
  wire  _T_1657 = _T_1656 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_182 = _T_1657 | _T_1666; // @[Reg.scala 28:19]
  wire  _T_1669 = _T_1652 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_1670 = _T_1651 & _T_1669; // @[Cache.scala 491:87]
  wire  _T_1671 = _T_1670 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_184 = _T_1671 | _T_1680; // @[Reg.scala 28:19]
  wire  _T_1683 = _T_1652 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_1684 = _T_1651 & _T_1683; // @[Cache.scala 491:87]
  wire  _T_1685 = _T_1684 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_186 = _T_1685 | _T_1694; // @[Reg.scala 28:19]
  wire  _T_1697 = _T_1652 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_1698 = _T_1651 & _T_1697; // @[Cache.scala 491:87]
  wire  _T_1699 = _T_1698 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_188 = _T_1699 | _T_1708; // @[Reg.scala 28:19]
  wire [1:0] _T_1710 = _T_1713 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_1712 = io_cacheOut_r_last_i & _T_189; // @[Cache.scala 488:28]
  wire  _T_1716 = _T_1713 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_1717 = _T_1712 & _T_1716; // @[Cache.scala 491:87]
  wire  _T_1718 = _T_1717 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_191 = _T_1718 | _T_1727; // @[Reg.scala 28:19]
  wire  _T_1730 = _T_1713 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_1731 = _T_1712 & _T_1730; // @[Cache.scala 491:87]
  wire  _T_1732 = _T_1731 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_193 = _T_1732 | _T_1741; // @[Reg.scala 28:19]
  wire  _T_1744 = _T_1713 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_1745 = _T_1712 & _T_1744; // @[Cache.scala 491:87]
  wire  _T_1746 = _T_1745 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_195 = _T_1746 | _T_1755; // @[Reg.scala 28:19]
  wire  _T_1758 = _T_1713 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_1759 = _T_1712 & _T_1758; // @[Cache.scala 491:87]
  wire  _T_1760 = _T_1759 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_197 = _T_1760 | _T_1769; // @[Reg.scala 28:19]
  wire [1:0] _T_1771 = _T_1774 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_1773 = io_cacheOut_r_last_i & _T_191; // @[Cache.scala 488:28]
  wire  _T_1777 = _T_1774 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_1778 = _T_1773 & _T_1777; // @[Cache.scala 491:87]
  wire  _T_1779 = _T_1778 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_200 = _T_1779 | _T_1788; // @[Reg.scala 28:19]
  wire  _T_1791 = _T_1774 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_1792 = _T_1773 & _T_1791; // @[Cache.scala 491:87]
  wire  _T_1793 = _T_1792 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_202 = _T_1793 | _T_1802; // @[Reg.scala 28:19]
  wire  _T_1805 = _T_1774 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_1806 = _T_1773 & _T_1805; // @[Cache.scala 491:87]
  wire  _T_1807 = _T_1806 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_204 = _T_1807 | _T_1816; // @[Reg.scala 28:19]
  wire  _T_1819 = _T_1774 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_1820 = _T_1773 & _T_1819; // @[Cache.scala 491:87]
  wire  _T_1821 = _T_1820 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_206 = _T_1821 | _T_1830; // @[Reg.scala 28:19]
  wire [1:0] _T_1832 = _T_1835 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_1834 = io_cacheOut_r_last_i & _T_193; // @[Cache.scala 488:28]
  wire  _T_1838 = _T_1835 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_1839 = _T_1834 & _T_1838; // @[Cache.scala 491:87]
  wire  _T_1840 = _T_1839 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_209 = _T_1840 | _T_1849; // @[Reg.scala 28:19]
  wire  _T_1852 = _T_1835 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_1853 = _T_1834 & _T_1852; // @[Cache.scala 491:87]
  wire  _T_1854 = _T_1853 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_211 = _T_1854 | _T_1863; // @[Reg.scala 28:19]
  wire  _T_1866 = _T_1835 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_1867 = _T_1834 & _T_1866; // @[Cache.scala 491:87]
  wire  _T_1868 = _T_1867 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_213 = _T_1868 | _T_1877; // @[Reg.scala 28:19]
  wire  _T_1880 = _T_1835 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_1881 = _T_1834 & _T_1880; // @[Cache.scala 491:87]
  wire  _T_1882 = _T_1881 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_215 = _T_1882 | _T_1891; // @[Reg.scala 28:19]
  wire [1:0] _T_1893 = _T_1896 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_1895 = io_cacheOut_r_last_i & _T_195; // @[Cache.scala 488:28]
  wire  _T_1899 = _T_1896 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_1900 = _T_1895 & _T_1899; // @[Cache.scala 491:87]
  wire  _T_1901 = _T_1900 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_218 = _T_1901 | _T_1910; // @[Reg.scala 28:19]
  wire  _T_1913 = _T_1896 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_1914 = _T_1895 & _T_1913; // @[Cache.scala 491:87]
  wire  _T_1915 = _T_1914 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_220 = _T_1915 | _T_1924; // @[Reg.scala 28:19]
  wire  _T_1927 = _T_1896 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_1928 = _T_1895 & _T_1927; // @[Cache.scala 491:87]
  wire  _T_1929 = _T_1928 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_222 = _T_1929 | _T_1938; // @[Reg.scala 28:19]
  wire  _T_1941 = _T_1896 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_1942 = _T_1895 & _T_1941; // @[Cache.scala 491:87]
  wire  _T_1943 = _T_1942 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_224 = _T_1943 | _T_1952; // @[Reg.scala 28:19]
  wire [1:0] _T_1954 = _T_1957 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_1956 = io_cacheOut_r_last_i & _T_197; // @[Cache.scala 488:28]
  wire  _T_1960 = _T_1957 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_1961 = _T_1956 & _T_1960; // @[Cache.scala 491:87]
  wire  _T_1962 = _T_1961 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_227 = _T_1962 | _T_1971; // @[Reg.scala 28:19]
  wire  _T_1974 = _T_1957 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_1975 = _T_1956 & _T_1974; // @[Cache.scala 491:87]
  wire  _T_1976 = _T_1975 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_229 = _T_1976 | _T_1985; // @[Reg.scala 28:19]
  wire  _T_1988 = _T_1957 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_1989 = _T_1956 & _T_1988; // @[Cache.scala 491:87]
  wire  _T_1990 = _T_1989 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_231 = _T_1990 | _T_1999; // @[Reg.scala 28:19]
  wire  _T_2002 = _T_1957 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_2003 = _T_1956 & _T_2002; // @[Cache.scala 491:87]
  wire  _T_2004 = _T_2003 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_233 = _T_2004 | _T_2013; // @[Reg.scala 28:19]
  wire [1:0] _T_2015 = _T_2018 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_2017 = io_cacheOut_r_last_i & _T_199; // @[Cache.scala 488:28]
  wire  _T_2021 = _T_2018 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_2022 = _T_2017 & _T_2021; // @[Cache.scala 491:87]
  wire  _T_2023 = _T_2022 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_236 = _T_2023 | _T_2032; // @[Reg.scala 28:19]
  wire  _T_2035 = _T_2018 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_2036 = _T_2017 & _T_2035; // @[Cache.scala 491:87]
  wire  _T_2037 = _T_2036 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_238 = _T_2037 | _T_2046; // @[Reg.scala 28:19]
  wire  _T_2049 = _T_2018 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_2050 = _T_2017 & _T_2049; // @[Cache.scala 491:87]
  wire  _T_2051 = _T_2050 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_240 = _T_2051 | _T_2060; // @[Reg.scala 28:19]
  wire  _T_2063 = _T_2018 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_2064 = _T_2017 & _T_2063; // @[Cache.scala 491:87]
  wire  _T_2065 = _T_2064 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_242 = _T_2065 | _T_2074; // @[Reg.scala 28:19]
  wire [1:0] _T_2076 = _T_2079 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_2078 = io_cacheOut_r_last_i & _T_201; // @[Cache.scala 488:28]
  wire  _T_2082 = _T_2079 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_2083 = _T_2078 & _T_2082; // @[Cache.scala 491:87]
  wire  _T_2084 = _T_2083 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_245 = _T_2084 | _T_2093; // @[Reg.scala 28:19]
  wire  _T_2096 = _T_2079 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_2097 = _T_2078 & _T_2096; // @[Cache.scala 491:87]
  wire  _T_2098 = _T_2097 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_247 = _T_2098 | _T_2107; // @[Reg.scala 28:19]
  wire  _T_2110 = _T_2079 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_2111 = _T_2078 & _T_2110; // @[Cache.scala 491:87]
  wire  _T_2112 = _T_2111 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_249 = _T_2112 | _T_2121; // @[Reg.scala 28:19]
  wire  _T_2124 = _T_2079 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_2125 = _T_2078 & _T_2124; // @[Cache.scala 491:87]
  wire  _T_2126 = _T_2125 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_251 = _T_2126 | _T_2135; // @[Reg.scala 28:19]
  wire [1:0] _T_2137 = _T_2140 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_2139 = io_cacheOut_r_last_i & _T_203; // @[Cache.scala 488:28]
  wire  _T_2143 = _T_2140 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_2144 = _T_2139 & _T_2143; // @[Cache.scala 491:87]
  wire  _T_2145 = _T_2144 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_254 = _T_2145 | _T_2154; // @[Reg.scala 28:19]
  wire  _T_2157 = _T_2140 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_2158 = _T_2139 & _T_2157; // @[Cache.scala 491:87]
  wire  _T_2159 = _T_2158 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_256 = _T_2159 | _T_2168; // @[Reg.scala 28:19]
  wire  _T_2171 = _T_2140 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_2172 = _T_2139 & _T_2171; // @[Cache.scala 491:87]
  wire  _T_2173 = _T_2172 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_258 = _T_2173 | _T_2182; // @[Reg.scala 28:19]
  wire  _T_2185 = _T_2140 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_2186 = _T_2139 & _T_2185; // @[Cache.scala 491:87]
  wire  _T_2187 = _T_2186 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_260 = _T_2187 | _T_2196; // @[Reg.scala 28:19]
  wire [1:0] _T_2198 = _T_2201 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_2200 = io_cacheOut_r_last_i & _T_205; // @[Cache.scala 488:28]
  wire  _T_2204 = _T_2201 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_2205 = _T_2200 & _T_2204; // @[Cache.scala 491:87]
  wire  _T_2206 = _T_2205 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_263 = _T_2206 | _T_2215; // @[Reg.scala 28:19]
  wire  _T_2218 = _T_2201 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_2219 = _T_2200 & _T_2218; // @[Cache.scala 491:87]
  wire  _T_2220 = _T_2219 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_265 = _T_2220 | _T_2229; // @[Reg.scala 28:19]
  wire  _T_2232 = _T_2201 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_2233 = _T_2200 & _T_2232; // @[Cache.scala 491:87]
  wire  _T_2234 = _T_2233 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_267 = _T_2234 | _T_2243; // @[Reg.scala 28:19]
  wire  _T_2246 = _T_2201 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_2247 = _T_2200 & _T_2246; // @[Cache.scala 491:87]
  wire  _T_2248 = _T_2247 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_269 = _T_2248 | _T_2257; // @[Reg.scala 28:19]
  wire [1:0] _T_2259 = _T_2262 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_2261 = io_cacheOut_r_last_i & _T_207; // @[Cache.scala 488:28]
  wire  _T_2265 = _T_2262 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_2266 = _T_2261 & _T_2265; // @[Cache.scala 491:87]
  wire  _T_2267 = _T_2266 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_272 = _T_2267 | _T_2276; // @[Reg.scala 28:19]
  wire  _T_2279 = _T_2262 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_2280 = _T_2261 & _T_2279; // @[Cache.scala 491:87]
  wire  _T_2281 = _T_2280 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_274 = _T_2281 | _T_2290; // @[Reg.scala 28:19]
  wire  _T_2293 = _T_2262 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_2294 = _T_2261 & _T_2293; // @[Cache.scala 491:87]
  wire  _T_2295 = _T_2294 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_276 = _T_2295 | _T_2304; // @[Reg.scala 28:19]
  wire  _T_2307 = _T_2262 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_2308 = _T_2261 & _T_2307; // @[Cache.scala 491:87]
  wire  _T_2309 = _T_2308 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_278 = _T_2309 | _T_2318; // @[Reg.scala 28:19]
  wire [1:0] _T_2320 = _T_2323 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_2322 = io_cacheOut_r_last_i & _T_209; // @[Cache.scala 488:28]
  wire  _T_2326 = _T_2323 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_2327 = _T_2322 & _T_2326; // @[Cache.scala 491:87]
  wire  _T_2328 = _T_2327 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_281 = _T_2328 | _T_2337; // @[Reg.scala 28:19]
  wire  _T_2340 = _T_2323 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_2341 = _T_2322 & _T_2340; // @[Cache.scala 491:87]
  wire  _T_2342 = _T_2341 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_283 = _T_2342 | _T_2351; // @[Reg.scala 28:19]
  wire  _T_2354 = _T_2323 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_2355 = _T_2322 & _T_2354; // @[Cache.scala 491:87]
  wire  _T_2356 = _T_2355 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_285 = _T_2356 | _T_2365; // @[Reg.scala 28:19]
  wire  _T_2368 = _T_2323 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_2369 = _T_2322 & _T_2368; // @[Cache.scala 491:87]
  wire  _T_2370 = _T_2369 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_287 = _T_2370 | _T_2379; // @[Reg.scala 28:19]
  wire [1:0] _T_2381 = _T_2384 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_2383 = io_cacheOut_r_last_i & _T_211; // @[Cache.scala 488:28]
  wire  _T_2387 = _T_2384 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_2388 = _T_2383 & _T_2387; // @[Cache.scala 491:87]
  wire  _T_2389 = _T_2388 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_290 = _T_2389 | _T_2398; // @[Reg.scala 28:19]
  wire  _T_2401 = _T_2384 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_2402 = _T_2383 & _T_2401; // @[Cache.scala 491:87]
  wire  _T_2403 = _T_2402 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_292 = _T_2403 | _T_2412; // @[Reg.scala 28:19]
  wire  _T_2415 = _T_2384 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_2416 = _T_2383 & _T_2415; // @[Cache.scala 491:87]
  wire  _T_2417 = _T_2416 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_294 = _T_2417 | _T_2426; // @[Reg.scala 28:19]
  wire  _T_2429 = _T_2384 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_2430 = _T_2383 & _T_2429; // @[Cache.scala 491:87]
  wire  _T_2431 = _T_2430 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_296 = _T_2431 | _T_2440; // @[Reg.scala 28:19]
  wire [1:0] _T_2442 = _T_2445 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_2444 = io_cacheOut_r_last_i & _T_213; // @[Cache.scala 488:28]
  wire  _T_2448 = _T_2445 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_2449 = _T_2444 & _T_2448; // @[Cache.scala 491:87]
  wire  _T_2450 = _T_2449 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_299 = _T_2450 | _T_2459; // @[Reg.scala 28:19]
  wire  _T_2462 = _T_2445 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_2463 = _T_2444 & _T_2462; // @[Cache.scala 491:87]
  wire  _T_2464 = _T_2463 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_301 = _T_2464 | _T_2473; // @[Reg.scala 28:19]
  wire  _T_2476 = _T_2445 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_2477 = _T_2444 & _T_2476; // @[Cache.scala 491:87]
  wire  _T_2478 = _T_2477 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_303 = _T_2478 | _T_2487; // @[Reg.scala 28:19]
  wire  _T_2490 = _T_2445 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_2491 = _T_2444 & _T_2490; // @[Cache.scala 491:87]
  wire  _T_2492 = _T_2491 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_305 = _T_2492 | _T_2501; // @[Reg.scala 28:19]
  wire [1:0] _T_2503 = _T_2506 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_2505 = io_cacheOut_r_last_i & _T_215; // @[Cache.scala 488:28]
  wire  _T_2509 = _T_2506 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_2510 = _T_2505 & _T_2509; // @[Cache.scala 491:87]
  wire  _T_2511 = _T_2510 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_308 = _T_2511 | _T_2520; // @[Reg.scala 28:19]
  wire  _T_2523 = _T_2506 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_2524 = _T_2505 & _T_2523; // @[Cache.scala 491:87]
  wire  _T_2525 = _T_2524 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_310 = _T_2525 | _T_2534; // @[Reg.scala 28:19]
  wire  _T_2537 = _T_2506 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_2538 = _T_2505 & _T_2537; // @[Cache.scala 491:87]
  wire  _T_2539 = _T_2538 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_312 = _T_2539 | _T_2548; // @[Reg.scala 28:19]
  wire  _T_2551 = _T_2506 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_2552 = _T_2505 & _T_2551; // @[Cache.scala 491:87]
  wire  _T_2553 = _T_2552 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_314 = _T_2553 | _T_2562; // @[Reg.scala 28:19]
  wire [1:0] _T_2564 = _T_2567 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_2566 = io_cacheOut_r_last_i & _T_217; // @[Cache.scala 488:28]
  wire  _T_2570 = _T_2567 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_2571 = _T_2566 & _T_2570; // @[Cache.scala 491:87]
  wire  _T_2572 = _T_2571 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_317 = _T_2572 | _T_2581; // @[Reg.scala 28:19]
  wire  _T_2584 = _T_2567 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_2585 = _T_2566 & _T_2584; // @[Cache.scala 491:87]
  wire  _T_2586 = _T_2585 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_319 = _T_2586 | _T_2595; // @[Reg.scala 28:19]
  wire  _T_2598 = _T_2567 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_2599 = _T_2566 & _T_2598; // @[Cache.scala 491:87]
  wire  _T_2600 = _T_2599 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_321 = _T_2600 | _T_2609; // @[Reg.scala 28:19]
  wire  _T_2612 = _T_2567 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_2613 = _T_2566 & _T_2612; // @[Cache.scala 491:87]
  wire  _T_2614 = _T_2613 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_323 = _T_2614 | _T_2623; // @[Reg.scala 28:19]
  wire [1:0] _T_2625 = _T_2628 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_2627 = io_cacheOut_r_last_i & _T_219; // @[Cache.scala 488:28]
  wire  _T_2631 = _T_2628 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_2632 = _T_2627 & _T_2631; // @[Cache.scala 491:87]
  wire  _T_2633 = _T_2632 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_326 = _T_2633 | _T_2642; // @[Reg.scala 28:19]
  wire  _T_2645 = _T_2628 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_2646 = _T_2627 & _T_2645; // @[Cache.scala 491:87]
  wire  _T_2647 = _T_2646 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_328 = _T_2647 | _T_2656; // @[Reg.scala 28:19]
  wire  _T_2659 = _T_2628 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_2660 = _T_2627 & _T_2659; // @[Cache.scala 491:87]
  wire  _T_2661 = _T_2660 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_330 = _T_2661 | _T_2670; // @[Reg.scala 28:19]
  wire  _T_2673 = _T_2628 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_2674 = _T_2627 & _T_2673; // @[Cache.scala 491:87]
  wire  _T_2675 = _T_2674 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_332 = _T_2675 | _T_2684; // @[Reg.scala 28:19]
  wire [1:0] _T_2686 = _T_2689 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_2688 = io_cacheOut_r_last_i & _T_221; // @[Cache.scala 488:28]
  wire  _T_2692 = _T_2689 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_2693 = _T_2688 & _T_2692; // @[Cache.scala 491:87]
  wire  _T_2694 = _T_2693 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_335 = _T_2694 | _T_2703; // @[Reg.scala 28:19]
  wire  _T_2706 = _T_2689 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_2707 = _T_2688 & _T_2706; // @[Cache.scala 491:87]
  wire  _T_2708 = _T_2707 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_337 = _T_2708 | _T_2717; // @[Reg.scala 28:19]
  wire  _T_2720 = _T_2689 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_2721 = _T_2688 & _T_2720; // @[Cache.scala 491:87]
  wire  _T_2722 = _T_2721 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_339 = _T_2722 | _T_2731; // @[Reg.scala 28:19]
  wire  _T_2734 = _T_2689 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_2735 = _T_2688 & _T_2734; // @[Cache.scala 491:87]
  wire  _T_2736 = _T_2735 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_341 = _T_2736 | _T_2745; // @[Reg.scala 28:19]
  wire [1:0] _T_2747 = _T_2750 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_2749 = io_cacheOut_r_last_i & _T_223; // @[Cache.scala 488:28]
  wire  _T_2753 = _T_2750 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_2754 = _T_2749 & _T_2753; // @[Cache.scala 491:87]
  wire  _T_2755 = _T_2754 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_344 = _T_2755 | _T_2764; // @[Reg.scala 28:19]
  wire  _T_2767 = _T_2750 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_2768 = _T_2749 & _T_2767; // @[Cache.scala 491:87]
  wire  _T_2769 = _T_2768 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_346 = _T_2769 | _T_2778; // @[Reg.scala 28:19]
  wire  _T_2781 = _T_2750 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_2782 = _T_2749 & _T_2781; // @[Cache.scala 491:87]
  wire  _T_2783 = _T_2782 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_348 = _T_2783 | _T_2792; // @[Reg.scala 28:19]
  wire  _T_2795 = _T_2750 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_2796 = _T_2749 & _T_2795; // @[Cache.scala 491:87]
  wire  _T_2797 = _T_2796 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_350 = _T_2797 | _T_2806; // @[Reg.scala 28:19]
  wire [1:0] _T_2808 = _T_2811 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_2810 = io_cacheOut_r_last_i & _T_225; // @[Cache.scala 488:28]
  wire  _T_2814 = _T_2811 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_2815 = _T_2810 & _T_2814; // @[Cache.scala 491:87]
  wire  _T_2816 = _T_2815 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_353 = _T_2816 | _T_2825; // @[Reg.scala 28:19]
  wire  _T_2828 = _T_2811 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_2829 = _T_2810 & _T_2828; // @[Cache.scala 491:87]
  wire  _T_2830 = _T_2829 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_355 = _T_2830 | _T_2839; // @[Reg.scala 28:19]
  wire  _T_2842 = _T_2811 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_2843 = _T_2810 & _T_2842; // @[Cache.scala 491:87]
  wire  _T_2844 = _T_2843 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_357 = _T_2844 | _T_2853; // @[Reg.scala 28:19]
  wire  _T_2856 = _T_2811 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_2857 = _T_2810 & _T_2856; // @[Cache.scala 491:87]
  wire  _T_2858 = _T_2857 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_359 = _T_2858 | _T_2867; // @[Reg.scala 28:19]
  wire [1:0] _T_2869 = _T_2872 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_2871 = io_cacheOut_r_last_i & _T_227; // @[Cache.scala 488:28]
  wire  _T_2875 = _T_2872 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_2876 = _T_2871 & _T_2875; // @[Cache.scala 491:87]
  wire  _T_2877 = _T_2876 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_362 = _T_2877 | _T_2886; // @[Reg.scala 28:19]
  wire  _T_2889 = _T_2872 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_2890 = _T_2871 & _T_2889; // @[Cache.scala 491:87]
  wire  _T_2891 = _T_2890 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_364 = _T_2891 | _T_2900; // @[Reg.scala 28:19]
  wire  _T_2903 = _T_2872 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_2904 = _T_2871 & _T_2903; // @[Cache.scala 491:87]
  wire  _T_2905 = _T_2904 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_366 = _T_2905 | _T_2914; // @[Reg.scala 28:19]
  wire  _T_2917 = _T_2872 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_2918 = _T_2871 & _T_2917; // @[Cache.scala 491:87]
  wire  _T_2919 = _T_2918 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_368 = _T_2919 | _T_2928; // @[Reg.scala 28:19]
  wire [1:0] _T_2930 = _T_2933 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_2932 = io_cacheOut_r_last_i & _T_229; // @[Cache.scala 488:28]
  wire  _T_2936 = _T_2933 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_2937 = _T_2932 & _T_2936; // @[Cache.scala 491:87]
  wire  _T_2938 = _T_2937 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_371 = _T_2938 | _T_2947; // @[Reg.scala 28:19]
  wire  _T_2950 = _T_2933 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_2951 = _T_2932 & _T_2950; // @[Cache.scala 491:87]
  wire  _T_2952 = _T_2951 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_373 = _T_2952 | _T_2961; // @[Reg.scala 28:19]
  wire  _T_2964 = _T_2933 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_2965 = _T_2932 & _T_2964; // @[Cache.scala 491:87]
  wire  _T_2966 = _T_2965 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_375 = _T_2966 | _T_2975; // @[Reg.scala 28:19]
  wire  _T_2978 = _T_2933 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_2979 = _T_2932 & _T_2978; // @[Cache.scala 491:87]
  wire  _T_2980 = _T_2979 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_377 = _T_2980 | _T_2989; // @[Reg.scala 28:19]
  wire [1:0] _T_2991 = _T_2994 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_2993 = io_cacheOut_r_last_i & _T_231; // @[Cache.scala 488:28]
  wire  _T_2997 = _T_2994 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_2998 = _T_2993 & _T_2997; // @[Cache.scala 491:87]
  wire  _T_2999 = _T_2998 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_380 = _T_2999 | _T_3008; // @[Reg.scala 28:19]
  wire  _T_3011 = _T_2994 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_3012 = _T_2993 & _T_3011; // @[Cache.scala 491:87]
  wire  _T_3013 = _T_3012 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_382 = _T_3013 | _T_3022; // @[Reg.scala 28:19]
  wire  _T_3025 = _T_2994 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_3026 = _T_2993 & _T_3025; // @[Cache.scala 491:87]
  wire  _T_3027 = _T_3026 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_384 = _T_3027 | _T_3036; // @[Reg.scala 28:19]
  wire  _T_3039 = _T_2994 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_3040 = _T_2993 & _T_3039; // @[Cache.scala 491:87]
  wire  _T_3041 = _T_3040 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_386 = _T_3041 | _T_3050; // @[Reg.scala 28:19]
  wire [1:0] _T_3052 = _T_3055 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_3054 = io_cacheOut_r_last_i & _T_233; // @[Cache.scala 488:28]
  wire  _T_3058 = _T_3055 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_3059 = _T_3054 & _T_3058; // @[Cache.scala 491:87]
  wire  _T_3060 = _T_3059 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_389 = _T_3060 | _T_3069; // @[Reg.scala 28:19]
  wire  _T_3072 = _T_3055 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_3073 = _T_3054 & _T_3072; // @[Cache.scala 491:87]
  wire  _T_3074 = _T_3073 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_391 = _T_3074 | _T_3083; // @[Reg.scala 28:19]
  wire  _T_3086 = _T_3055 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_3087 = _T_3054 & _T_3086; // @[Cache.scala 491:87]
  wire  _T_3088 = _T_3087 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_393 = _T_3088 | _T_3097; // @[Reg.scala 28:19]
  wire  _T_3100 = _T_3055 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_3101 = _T_3054 & _T_3100; // @[Cache.scala 491:87]
  wire  _T_3102 = _T_3101 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_395 = _T_3102 | _T_3111; // @[Reg.scala 28:19]
  wire [1:0] _T_3113 = _T_3116 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_3115 = io_cacheOut_r_last_i & _T_235; // @[Cache.scala 488:28]
  wire  _T_3119 = _T_3116 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_3120 = _T_3115 & _T_3119; // @[Cache.scala 491:87]
  wire  _T_3121 = _T_3120 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_398 = _T_3121 | _T_3130; // @[Reg.scala 28:19]
  wire  _T_3133 = _T_3116 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_3134 = _T_3115 & _T_3133; // @[Cache.scala 491:87]
  wire  _T_3135 = _T_3134 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_400 = _T_3135 | _T_3144; // @[Reg.scala 28:19]
  wire  _T_3147 = _T_3116 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_3148 = _T_3115 & _T_3147; // @[Cache.scala 491:87]
  wire  _T_3149 = _T_3148 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_402 = _T_3149 | _T_3158; // @[Reg.scala 28:19]
  wire  _T_3161 = _T_3116 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_3162 = _T_3115 & _T_3161; // @[Cache.scala 491:87]
  wire  _T_3163 = _T_3162 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_404 = _T_3163 | _T_3172; // @[Reg.scala 28:19]
  wire [1:0] _T_3174 = _T_3177 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_3176 = io_cacheOut_r_last_i & _T_237; // @[Cache.scala 488:28]
  wire  _T_3180 = _T_3177 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_3181 = _T_3176 & _T_3180; // @[Cache.scala 491:87]
  wire  _T_3182 = _T_3181 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_407 = _T_3182 | _T_3191; // @[Reg.scala 28:19]
  wire  _T_3194 = _T_3177 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_3195 = _T_3176 & _T_3194; // @[Cache.scala 491:87]
  wire  _T_3196 = _T_3195 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_409 = _T_3196 | _T_3205; // @[Reg.scala 28:19]
  wire  _T_3208 = _T_3177 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_3209 = _T_3176 & _T_3208; // @[Cache.scala 491:87]
  wire  _T_3210 = _T_3209 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_411 = _T_3210 | _T_3219; // @[Reg.scala 28:19]
  wire  _T_3222 = _T_3177 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_3223 = _T_3176 & _T_3222; // @[Cache.scala 491:87]
  wire  _T_3224 = _T_3223 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_413 = _T_3224 | _T_3233; // @[Reg.scala 28:19]
  wire [1:0] _T_3235 = _T_3238 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_3237 = io_cacheOut_r_last_i & _T_239; // @[Cache.scala 488:28]
  wire  _T_3241 = _T_3238 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_3242 = _T_3237 & _T_3241; // @[Cache.scala 491:87]
  wire  _T_3243 = _T_3242 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_416 = _T_3243 | _T_3252; // @[Reg.scala 28:19]
  wire  _T_3255 = _T_3238 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_3256 = _T_3237 & _T_3255; // @[Cache.scala 491:87]
  wire  _T_3257 = _T_3256 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_418 = _T_3257 | _T_3266; // @[Reg.scala 28:19]
  wire  _T_3269 = _T_3238 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_3270 = _T_3237 & _T_3269; // @[Cache.scala 491:87]
  wire  _T_3271 = _T_3270 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_420 = _T_3271 | _T_3280; // @[Reg.scala 28:19]
  wire  _T_3283 = _T_3238 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_3284 = _T_3237 & _T_3283; // @[Cache.scala 491:87]
  wire  _T_3285 = _T_3284 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_422 = _T_3285 | _T_3294; // @[Reg.scala 28:19]
  wire [1:0] _T_3296 = _T_3299 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_3298 = io_cacheOut_r_last_i & _T_241; // @[Cache.scala 488:28]
  wire  _T_3302 = _T_3299 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_3303 = _T_3298 & _T_3302; // @[Cache.scala 491:87]
  wire  _T_3304 = _T_3303 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_425 = _T_3304 | _T_3313; // @[Reg.scala 28:19]
  wire  _T_3316 = _T_3299 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_3317 = _T_3298 & _T_3316; // @[Cache.scala 491:87]
  wire  _T_3318 = _T_3317 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_427 = _T_3318 | _T_3327; // @[Reg.scala 28:19]
  wire  _T_3330 = _T_3299 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_3331 = _T_3298 & _T_3330; // @[Cache.scala 491:87]
  wire  _T_3332 = _T_3331 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_429 = _T_3332 | _T_3341; // @[Reg.scala 28:19]
  wire  _T_3344 = _T_3299 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_3345 = _T_3298 & _T_3344; // @[Cache.scala 491:87]
  wire  _T_3346 = _T_3345 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_431 = _T_3346 | _T_3355; // @[Reg.scala 28:19]
  wire [1:0] _T_3357 = _T_3360 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_3359 = io_cacheOut_r_last_i & _T_243; // @[Cache.scala 488:28]
  wire  _T_3363 = _T_3360 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_3364 = _T_3359 & _T_3363; // @[Cache.scala 491:87]
  wire  _T_3365 = _T_3364 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_434 = _T_3365 | _T_3374; // @[Reg.scala 28:19]
  wire  _T_3377 = _T_3360 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_3378 = _T_3359 & _T_3377; // @[Cache.scala 491:87]
  wire  _T_3379 = _T_3378 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_436 = _T_3379 | _T_3388; // @[Reg.scala 28:19]
  wire  _T_3391 = _T_3360 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_3392 = _T_3359 & _T_3391; // @[Cache.scala 491:87]
  wire  _T_3393 = _T_3392 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_438 = _T_3393 | _T_3402; // @[Reg.scala 28:19]
  wire  _T_3405 = _T_3360 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_3406 = _T_3359 & _T_3405; // @[Cache.scala 491:87]
  wire  _T_3407 = _T_3406 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_440 = _T_3407 | _T_3416; // @[Reg.scala 28:19]
  wire [1:0] _T_3418 = _T_3421 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_3420 = io_cacheOut_r_last_i & _T_245; // @[Cache.scala 488:28]
  wire  _T_3424 = _T_3421 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_3425 = _T_3420 & _T_3424; // @[Cache.scala 491:87]
  wire  _T_3426 = _T_3425 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_443 = _T_3426 | _T_3435; // @[Reg.scala 28:19]
  wire  _T_3438 = _T_3421 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_3439 = _T_3420 & _T_3438; // @[Cache.scala 491:87]
  wire  _T_3440 = _T_3439 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_445 = _T_3440 | _T_3449; // @[Reg.scala 28:19]
  wire  _T_3452 = _T_3421 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_3453 = _T_3420 & _T_3452; // @[Cache.scala 491:87]
  wire  _T_3454 = _T_3453 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_447 = _T_3454 | _T_3463; // @[Reg.scala 28:19]
  wire  _T_3466 = _T_3421 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_3467 = _T_3420 & _T_3466; // @[Cache.scala 491:87]
  wire  _T_3468 = _T_3467 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_449 = _T_3468 | _T_3477; // @[Reg.scala 28:19]
  wire [1:0] _T_3479 = _T_3482 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_3481 = io_cacheOut_r_last_i & _T_247; // @[Cache.scala 488:28]
  wire  _T_3485 = _T_3482 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_3486 = _T_3481 & _T_3485; // @[Cache.scala 491:87]
  wire  _T_3487 = _T_3486 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_452 = _T_3487 | _T_3496; // @[Reg.scala 28:19]
  wire  _T_3499 = _T_3482 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_3500 = _T_3481 & _T_3499; // @[Cache.scala 491:87]
  wire  _T_3501 = _T_3500 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_454 = _T_3501 | _T_3510; // @[Reg.scala 28:19]
  wire  _T_3513 = _T_3482 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_3514 = _T_3481 & _T_3513; // @[Cache.scala 491:87]
  wire  _T_3515 = _T_3514 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_456 = _T_3515 | _T_3524; // @[Reg.scala 28:19]
  wire  _T_3527 = _T_3482 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_3528 = _T_3481 & _T_3527; // @[Cache.scala 491:87]
  wire  _T_3529 = _T_3528 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_458 = _T_3529 | _T_3538; // @[Reg.scala 28:19]
  wire [1:0] _T_3540 = _T_3543 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_3542 = io_cacheOut_r_last_i & _T_249; // @[Cache.scala 488:28]
  wire  _T_3546 = _T_3543 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_3547 = _T_3542 & _T_3546; // @[Cache.scala 491:87]
  wire  _T_3548 = _T_3547 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_461 = _T_3548 | _T_3557; // @[Reg.scala 28:19]
  wire  _T_3560 = _T_3543 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_3561 = _T_3542 & _T_3560; // @[Cache.scala 491:87]
  wire  _T_3562 = _T_3561 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_463 = _T_3562 | _T_3571; // @[Reg.scala 28:19]
  wire  _T_3574 = _T_3543 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_3575 = _T_3542 & _T_3574; // @[Cache.scala 491:87]
  wire  _T_3576 = _T_3575 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_465 = _T_3576 | _T_3585; // @[Reg.scala 28:19]
  wire  _T_3588 = _T_3543 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_3589 = _T_3542 & _T_3588; // @[Cache.scala 491:87]
  wire  _T_3590 = _T_3589 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_467 = _T_3590 | _T_3599; // @[Reg.scala 28:19]
  wire [1:0] _T_3601 = _T_3604 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_3603 = io_cacheOut_r_last_i & _T_251; // @[Cache.scala 488:28]
  wire  _T_3607 = _T_3604 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_3608 = _T_3603 & _T_3607; // @[Cache.scala 491:87]
  wire  _T_3609 = _T_3608 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_470 = _T_3609 | _T_3618; // @[Reg.scala 28:19]
  wire  _T_3621 = _T_3604 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_3622 = _T_3603 & _T_3621; // @[Cache.scala 491:87]
  wire  _T_3623 = _T_3622 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_472 = _T_3623 | _T_3632; // @[Reg.scala 28:19]
  wire  _T_3635 = _T_3604 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_3636 = _T_3603 & _T_3635; // @[Cache.scala 491:87]
  wire  _T_3637 = _T_3636 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_474 = _T_3637 | _T_3646; // @[Reg.scala 28:19]
  wire  _T_3649 = _T_3604 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_3650 = _T_3603 & _T_3649; // @[Cache.scala 491:87]
  wire  _T_3651 = _T_3650 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_476 = _T_3651 | _T_3660; // @[Reg.scala 28:19]
  wire [1:0] _T_3662 = _T_3665 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_3664 = io_cacheOut_r_last_i & _T_253; // @[Cache.scala 488:28]
  wire  _T_3668 = _T_3665 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_3669 = _T_3664 & _T_3668; // @[Cache.scala 491:87]
  wire  _T_3670 = _T_3669 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_479 = _T_3670 | _T_3679; // @[Reg.scala 28:19]
  wire  _T_3682 = _T_3665 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_3683 = _T_3664 & _T_3682; // @[Cache.scala 491:87]
  wire  _T_3684 = _T_3683 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_481 = _T_3684 | _T_3693; // @[Reg.scala 28:19]
  wire  _T_3696 = _T_3665 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_3697 = _T_3664 & _T_3696; // @[Cache.scala 491:87]
  wire  _T_3698 = _T_3697 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_483 = _T_3698 | _T_3707; // @[Reg.scala 28:19]
  wire  _T_3710 = _T_3665 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_3711 = _T_3664 & _T_3710; // @[Cache.scala 491:87]
  wire  _T_3712 = _T_3711 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_485 = _T_3712 | _T_3721; // @[Reg.scala 28:19]
  wire [1:0] _T_3723 = _T_3726 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_3725 = io_cacheOut_r_last_i & _T_255; // @[Cache.scala 488:28]
  wire  _T_3729 = _T_3726 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_3730 = _T_3725 & _T_3729; // @[Cache.scala 491:87]
  wire  _T_3731 = _T_3730 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_488 = _T_3731 | _T_3740; // @[Reg.scala 28:19]
  wire  _T_3743 = _T_3726 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_3744 = _T_3725 & _T_3743; // @[Cache.scala 491:87]
  wire  _T_3745 = _T_3744 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_490 = _T_3745 | _T_3754; // @[Reg.scala 28:19]
  wire  _T_3757 = _T_3726 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_3758 = _T_3725 & _T_3757; // @[Cache.scala 491:87]
  wire  _T_3759 = _T_3758 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_492 = _T_3759 | _T_3768; // @[Reg.scala 28:19]
  wire  _T_3771 = _T_3726 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_3772 = _T_3725 & _T_3771; // @[Cache.scala 491:87]
  wire  _T_3773 = _T_3772 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_494 = _T_3773 | _T_3782; // @[Reg.scala 28:19]
  wire [1:0] _T_3784 = _T_3787 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_3786 = io_cacheOut_r_last_i & _T_257; // @[Cache.scala 488:28]
  wire  _T_3790 = _T_3787 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_3791 = _T_3786 & _T_3790; // @[Cache.scala 491:87]
  wire  _T_3792 = _T_3791 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_497 = _T_3792 | _T_3801; // @[Reg.scala 28:19]
  wire  _T_3804 = _T_3787 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_3805 = _T_3786 & _T_3804; // @[Cache.scala 491:87]
  wire  _T_3806 = _T_3805 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_499 = _T_3806 | _T_3815; // @[Reg.scala 28:19]
  wire  _T_3818 = _T_3787 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_3819 = _T_3786 & _T_3818; // @[Cache.scala 491:87]
  wire  _T_3820 = _T_3819 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_501 = _T_3820 | _T_3829; // @[Reg.scala 28:19]
  wire  _T_3832 = _T_3787 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_3833 = _T_3786 & _T_3832; // @[Cache.scala 491:87]
  wire  _T_3834 = _T_3833 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_503 = _T_3834 | _T_3843; // @[Reg.scala 28:19]
  wire [1:0] _T_3845 = _T_3848 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_3847 = io_cacheOut_r_last_i & _T_259; // @[Cache.scala 488:28]
  wire  _T_3851 = _T_3848 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_3852 = _T_3847 & _T_3851; // @[Cache.scala 491:87]
  wire  _T_3853 = _T_3852 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_506 = _T_3853 | _T_3862; // @[Reg.scala 28:19]
  wire  _T_3865 = _T_3848 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_3866 = _T_3847 & _T_3865; // @[Cache.scala 491:87]
  wire  _T_3867 = _T_3866 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_508 = _T_3867 | _T_3876; // @[Reg.scala 28:19]
  wire  _T_3879 = _T_3848 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_3880 = _T_3847 & _T_3879; // @[Cache.scala 491:87]
  wire  _T_3881 = _T_3880 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_510 = _T_3881 | _T_3890; // @[Reg.scala 28:19]
  wire  _T_3893 = _T_3848 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_3894 = _T_3847 & _T_3893; // @[Cache.scala 491:87]
  wire  _T_3895 = _T_3894 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_512 = _T_3895 | _T_3904; // @[Reg.scala 28:19]
  wire [1:0] _T_3906 = _T_3909 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_3908 = io_cacheOut_r_last_i & _T_261; // @[Cache.scala 488:28]
  wire  _T_3912 = _T_3909 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_3913 = _T_3908 & _T_3912; // @[Cache.scala 491:87]
  wire  _T_3914 = _T_3913 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_515 = _T_3914 | _T_3923; // @[Reg.scala 28:19]
  wire  _T_3926 = _T_3909 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_3927 = _T_3908 & _T_3926; // @[Cache.scala 491:87]
  wire  _T_3928 = _T_3927 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_517 = _T_3928 | _T_3937; // @[Reg.scala 28:19]
  wire  _T_3940 = _T_3909 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_3941 = _T_3908 & _T_3940; // @[Cache.scala 491:87]
  wire  _T_3942 = _T_3941 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_519 = _T_3942 | _T_3951; // @[Reg.scala 28:19]
  wire  _T_3954 = _T_3909 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_3955 = _T_3908 & _T_3954; // @[Cache.scala 491:87]
  wire  _T_3956 = _T_3955 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_521 = _T_3956 | _T_3965; // @[Reg.scala 28:19]
  wire [1:0] _T_3967 = _T_3970 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_3969 = io_cacheOut_r_last_i & _T_263; // @[Cache.scala 488:28]
  wire  _T_3973 = _T_3970 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_3974 = _T_3969 & _T_3973; // @[Cache.scala 491:87]
  wire  _T_3975 = _T_3974 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_524 = _T_3975 | _T_3984; // @[Reg.scala 28:19]
  wire  _T_3987 = _T_3970 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_3988 = _T_3969 & _T_3987; // @[Cache.scala 491:87]
  wire  _T_3989 = _T_3988 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_526 = _T_3989 | _T_3998; // @[Reg.scala 28:19]
  wire  _T_4001 = _T_3970 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_4002 = _T_3969 & _T_4001; // @[Cache.scala 491:87]
  wire  _T_4003 = _T_4002 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_528 = _T_4003 | _T_4012; // @[Reg.scala 28:19]
  wire  _T_4015 = _T_3970 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_4016 = _T_3969 & _T_4015; // @[Cache.scala 491:87]
  wire  _T_4017 = _T_4016 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_530 = _T_4017 | _T_4026; // @[Reg.scala 28:19]
  wire [1:0] _T_4028 = _T_4031 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_4030 = io_cacheOut_r_last_i & _T_265; // @[Cache.scala 488:28]
  wire  _T_4034 = _T_4031 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_4035 = _T_4030 & _T_4034; // @[Cache.scala 491:87]
  wire  _T_4036 = _T_4035 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_533 = _T_4036 | _T_4045; // @[Reg.scala 28:19]
  wire  _T_4048 = _T_4031 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_4049 = _T_4030 & _T_4048; // @[Cache.scala 491:87]
  wire  _T_4050 = _T_4049 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_535 = _T_4050 | _T_4059; // @[Reg.scala 28:19]
  wire  _T_4062 = _T_4031 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_4063 = _T_4030 & _T_4062; // @[Cache.scala 491:87]
  wire  _T_4064 = _T_4063 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_537 = _T_4064 | _T_4073; // @[Reg.scala 28:19]
  wire  _T_4076 = _T_4031 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_4077 = _T_4030 & _T_4076; // @[Cache.scala 491:87]
  wire  _T_4078 = _T_4077 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_539 = _T_4078 | _T_4087; // @[Reg.scala 28:19]
  wire [1:0] _T_4089 = _T_4092 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_4091 = io_cacheOut_r_last_i & _T_267; // @[Cache.scala 488:28]
  wire  _T_4095 = _T_4092 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_4096 = _T_4091 & _T_4095; // @[Cache.scala 491:87]
  wire  _T_4097 = _T_4096 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_542 = _T_4097 | _T_4106; // @[Reg.scala 28:19]
  wire  _T_4109 = _T_4092 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_4110 = _T_4091 & _T_4109; // @[Cache.scala 491:87]
  wire  _T_4111 = _T_4110 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_544 = _T_4111 | _T_4120; // @[Reg.scala 28:19]
  wire  _T_4123 = _T_4092 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_4124 = _T_4091 & _T_4123; // @[Cache.scala 491:87]
  wire  _T_4125 = _T_4124 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_546 = _T_4125 | _T_4134; // @[Reg.scala 28:19]
  wire  _T_4137 = _T_4092 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_4138 = _T_4091 & _T_4137; // @[Cache.scala 491:87]
  wire  _T_4139 = _T_4138 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_548 = _T_4139 | _T_4148; // @[Reg.scala 28:19]
  wire [1:0] _T_4150 = _T_4153 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_4152 = io_cacheOut_r_last_i & _T_269; // @[Cache.scala 488:28]
  wire  _T_4156 = _T_4153 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_4157 = _T_4152 & _T_4156; // @[Cache.scala 491:87]
  wire  _T_4158 = _T_4157 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_551 = _T_4158 | _T_4167; // @[Reg.scala 28:19]
  wire  _T_4170 = _T_4153 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_4171 = _T_4152 & _T_4170; // @[Cache.scala 491:87]
  wire  _T_4172 = _T_4171 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_553 = _T_4172 | _T_4181; // @[Reg.scala 28:19]
  wire  _T_4184 = _T_4153 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_4185 = _T_4152 & _T_4184; // @[Cache.scala 491:87]
  wire  _T_4186 = _T_4185 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_555 = _T_4186 | _T_4195; // @[Reg.scala 28:19]
  wire  _T_4198 = _T_4153 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_4199 = _T_4152 & _T_4198; // @[Cache.scala 491:87]
  wire  _T_4200 = _T_4199 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_557 = _T_4200 | _T_4209; // @[Reg.scala 28:19]
  wire [1:0] _T_4211 = _T_4214 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_4213 = io_cacheOut_r_last_i & _T_271; // @[Cache.scala 488:28]
  wire  _T_4217 = _T_4214 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_4218 = _T_4213 & _T_4217; // @[Cache.scala 491:87]
  wire  _T_4219 = _T_4218 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_560 = _T_4219 | _T_4228; // @[Reg.scala 28:19]
  wire  _T_4231 = _T_4214 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_4232 = _T_4213 & _T_4231; // @[Cache.scala 491:87]
  wire  _T_4233 = _T_4232 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_562 = _T_4233 | _T_4242; // @[Reg.scala 28:19]
  wire  _T_4245 = _T_4214 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_4246 = _T_4213 & _T_4245; // @[Cache.scala 491:87]
  wire  _T_4247 = _T_4246 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_564 = _T_4247 | _T_4256; // @[Reg.scala 28:19]
  wire  _T_4259 = _T_4214 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_4260 = _T_4213 & _T_4259; // @[Cache.scala 491:87]
  wire  _T_4261 = _T_4260 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_566 = _T_4261 | _T_4270; // @[Reg.scala 28:19]
  wire [1:0] _T_4272 = _T_4275 + 2'h1; // @[Cache.scala 486:23]
  wire  _T_4274 = io_cacheOut_r_last_i & _T_273; // @[Cache.scala 488:28]
  wire  _T_4278 = _T_4275 == 2'h0; // @[Cache.scala 491:106]
  wire  _T_4279 = _T_4274 & _T_4278; // @[Cache.scala 491:87]
  wire  _T_4280 = _T_4279 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_569 = _T_4280 | _T_4289; // @[Reg.scala 28:19]
  wire  _T_4292 = _T_4275 == 2'h1; // @[Cache.scala 491:106]
  wire  _T_4293 = _T_4274 & _T_4292; // @[Cache.scala 491:87]
  wire  _T_4294 = _T_4293 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_571 = _T_4294 | _T_4303; // @[Reg.scala 28:19]
  wire  _T_4306 = _T_4275 == 2'h2; // @[Cache.scala 491:106]
  wire  _T_4307 = _T_4274 & _T_4306; // @[Cache.scala 491:87]
  wire  _T_4308 = _T_4307 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_573 = _T_4308 | _T_4317; // @[Reg.scala 28:19]
  wire  _T_4320 = _T_4275 == 2'h3; // @[Cache.scala 491:106]
  wire  _T_4321 = _T_4274 & _T_4320; // @[Cache.scala 491:87]
  wire  _T_4322 = _T_4321 & _T_18; // @[Cache.scala 491:114]
  wire  _GEN_575 = _T_4322 | _T_4331; // @[Reg.scala 28:19]
  wire  _T_4387 = _T_18 & io_cacheOut_r_valid_i; // @[Cache.scala 524:27]
  wire  _T_4388 = 2'h0 == _T_425; // @[Cache.scala 524:62]
  wire  _T_4389 = _T_4387 & _T_4388; // @[Cache.scala 524:53]
  wire  _T_4390 = io_cacheIn_valid & _T_276; // @[Cache.scala 524:96]
  wire  _T_4391 = _T_4390 & _T_17; // @[Cache.scala 524:113]
  wire  _T_4392 = _T_4389 | _T_4391; // @[Cache.scala 524:75]
  wire [127:0] _T_4400 = {io_cacheOut_r_data_i,64'h0}; // @[Cat.scala 29:58]
  wire [127:0] _T_4401 = {64'h0,io_cacheOut_r_data_i}; // @[Cat.scala 29:58]
  wire  _T_4411 = 2'h1 == _T_425; // @[Cache.scala 524:62]
  wire  _T_4412 = _T_4387 & _T_4411; // @[Cache.scala 524:53]
  wire  _T_4413 = io_cacheIn_valid & _T_278; // @[Cache.scala 524:96]
  wire  _T_4414 = _T_4413 & _T_17; // @[Cache.scala 524:113]
  wire  _T_4415 = _T_4412 | _T_4414; // @[Cache.scala 524:75]
  wire  _T_4434 = 2'h2 == _T_425; // @[Cache.scala 524:62]
  wire  _T_4435 = _T_4387 & _T_4434; // @[Cache.scala 524:53]
  wire  _T_4436 = io_cacheIn_valid & _T_280; // @[Cache.scala 524:96]
  wire  _T_4437 = _T_4436 & _T_17; // @[Cache.scala 524:113]
  wire  _T_4438 = _T_4435 | _T_4437; // @[Cache.scala 524:75]
  wire  _T_4457 = 2'h3 == _T_425; // @[Cache.scala 524:62]
  wire  _T_4458 = _T_4387 & _T_4457; // @[Cache.scala 524:53]
  wire  _T_4459 = io_cacheIn_valid & _T_282; // @[Cache.scala 524:96]
  wire  _T_4460 = _T_4459 & _T_17; // @[Cache.scala 524:113]
  wire  _T_4461 = _T_4458 | _T_4460; // @[Cache.scala 524:75]
  assign io_cacheOut_ar_valid_o = _T_4 == 2'h1; // @[Cache.scala 482:26]
  assign io_cacheOut_ar_addr_o = {io_cacheIn_addr[31:4],4'h0}; // @[Cache.scala 481:25]
  assign io_cacheOut_ar_len_o = {{7'd0}, _T_18}; // @[Cache.scala 480:24]
  assign io_cacheOut_w_addr_o = io_cacheIn_addr; // @[Cache.scala 516:24]
  assign io_cacheIn_ready = _T_19 | _T_20; // @[Cache.scala 532:20]
  assign io_cacheIn_data_read = io_cacheIn_addr[3] ? _T_293[127:64] : _T_293[63:0]; // @[Cache.scala 466:24]
  assign io_SRAMIO_0_cen = ~_T_4392; // @[Cache.scala 524:13]
  assign io_SRAMIO_0_wen = ~_T_4389; // @[Cache.scala 526:13]
  assign io_SRAMIO_0_wdata = io_cacheOut_r_last_i ? _T_4400 : _T_4401; // @[Cache.scala 527:15]
  assign io_SRAMIO_0_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 525:14]
  assign io_SRAMIO_0_wmask = io_cacheOut_r_last_i ? 128'hffffffffffffffff : 128'hffffffffffffffff0000000000000000; // @[Cache.scala 528:15]
  assign io_SRAMIO_1_cen = ~_T_4415; // @[Cache.scala 524:13]
  assign io_SRAMIO_1_wen = ~_T_4412; // @[Cache.scala 526:13]
  assign io_SRAMIO_1_wdata = io_cacheOut_r_last_i ? _T_4400 : _T_4401; // @[Cache.scala 527:15]
  assign io_SRAMIO_1_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 525:14]
  assign io_SRAMIO_1_wmask = io_cacheOut_r_last_i ? 128'hffffffffffffffff : 128'hffffffffffffffff0000000000000000; // @[Cache.scala 528:15]
  assign io_SRAMIO_2_cen = ~_T_4438; // @[Cache.scala 524:13]
  assign io_SRAMIO_2_wen = ~_T_4435; // @[Cache.scala 526:13]
  assign io_SRAMIO_2_wdata = io_cacheOut_r_last_i ? _T_4400 : _T_4401; // @[Cache.scala 527:15]
  assign io_SRAMIO_2_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 525:14]
  assign io_SRAMIO_2_wmask = io_cacheOut_r_last_i ? 128'hffffffffffffffff : 128'hffffffffffffffff0000000000000000; // @[Cache.scala 528:15]
  assign io_SRAMIO_3_cen = ~_T_4461; // @[Cache.scala 524:13]
  assign io_SRAMIO_3_wen = ~_T_4458; // @[Cache.scala 526:13]
  assign io_SRAMIO_3_wdata = io_cacheOut_r_last_i ? _T_4400 : _T_4401; // @[Cache.scala 527:15]
  assign io_SRAMIO_3_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 525:14]
  assign io_SRAMIO_3_wmask = io_cacheOut_r_last_i ? 128'hffffffffffffffff : 128'hffffffffffffffff0000000000000000; // @[Cache.scala 528:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_4 = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  _T_4289 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_4228 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _T_4167 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_4106 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_4045 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_3984 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_3923 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_3862 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_3801 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_3740 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_3679 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_3618 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_3557 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_3496 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_3435 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _T_3374 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _T_3313 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_3252 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _T_3191 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _T_3130 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_3069 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  _T_3008 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _T_2947 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  _T_2886 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  _T_2825 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  _T_2764 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  _T_2703 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  _T_2642 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  _T_2581 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  _T_2520 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  _T_2459 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  _T_2398 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  _T_2337 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  _T_2276 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  _T_2215 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  _T_2154 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  _T_2093 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  _T_2032 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  _T_1971 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  _T_1910 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  _T_1849 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  _T_1788 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  _T_1727 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  _T_1666 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  _T_1605 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  _T_1544 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  _T_1483 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  _T_1422 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  _T_1361 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  _T_1300 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  _T_1239 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  _T_1178 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  _T_1117 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  _T_1056 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  _T_995 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  _T_934 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  _T_873 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  _T_812 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  _T_751 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  _T_690 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  _T_629 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  _T_568 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  _T_507 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  _T_446 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  _T_4281 = _RAND_65[21:0];
  _RAND_66 = {1{`RANDOM}};
  _T_4220 = _RAND_66[21:0];
  _RAND_67 = {1{`RANDOM}};
  _T_4159 = _RAND_67[21:0];
  _RAND_68 = {1{`RANDOM}};
  _T_4098 = _RAND_68[21:0];
  _RAND_69 = {1{`RANDOM}};
  _T_4037 = _RAND_69[21:0];
  _RAND_70 = {1{`RANDOM}};
  _T_3976 = _RAND_70[21:0];
  _RAND_71 = {1{`RANDOM}};
  _T_3915 = _RAND_71[21:0];
  _RAND_72 = {1{`RANDOM}};
  _T_3854 = _RAND_72[21:0];
  _RAND_73 = {1{`RANDOM}};
  _T_3793 = _RAND_73[21:0];
  _RAND_74 = {1{`RANDOM}};
  _T_3732 = _RAND_74[21:0];
  _RAND_75 = {1{`RANDOM}};
  _T_3671 = _RAND_75[21:0];
  _RAND_76 = {1{`RANDOM}};
  _T_3610 = _RAND_76[21:0];
  _RAND_77 = {1{`RANDOM}};
  _T_3549 = _RAND_77[21:0];
  _RAND_78 = {1{`RANDOM}};
  _T_3488 = _RAND_78[21:0];
  _RAND_79 = {1{`RANDOM}};
  _T_3427 = _RAND_79[21:0];
  _RAND_80 = {1{`RANDOM}};
  _T_3366 = _RAND_80[21:0];
  _RAND_81 = {1{`RANDOM}};
  _T_3305 = _RAND_81[21:0];
  _RAND_82 = {1{`RANDOM}};
  _T_3244 = _RAND_82[21:0];
  _RAND_83 = {1{`RANDOM}};
  _T_3183 = _RAND_83[21:0];
  _RAND_84 = {1{`RANDOM}};
  _T_3122 = _RAND_84[21:0];
  _RAND_85 = {1{`RANDOM}};
  _T_3061 = _RAND_85[21:0];
  _RAND_86 = {1{`RANDOM}};
  _T_3000 = _RAND_86[21:0];
  _RAND_87 = {1{`RANDOM}};
  _T_2939 = _RAND_87[21:0];
  _RAND_88 = {1{`RANDOM}};
  _T_2878 = _RAND_88[21:0];
  _RAND_89 = {1{`RANDOM}};
  _T_2817 = _RAND_89[21:0];
  _RAND_90 = {1{`RANDOM}};
  _T_2756 = _RAND_90[21:0];
  _RAND_91 = {1{`RANDOM}};
  _T_2695 = _RAND_91[21:0];
  _RAND_92 = {1{`RANDOM}};
  _T_2634 = _RAND_92[21:0];
  _RAND_93 = {1{`RANDOM}};
  _T_2573 = _RAND_93[21:0];
  _RAND_94 = {1{`RANDOM}};
  _T_2512 = _RAND_94[21:0];
  _RAND_95 = {1{`RANDOM}};
  _T_2451 = _RAND_95[21:0];
  _RAND_96 = {1{`RANDOM}};
  _T_2390 = _RAND_96[21:0];
  _RAND_97 = {1{`RANDOM}};
  _T_2329 = _RAND_97[21:0];
  _RAND_98 = {1{`RANDOM}};
  _T_2268 = _RAND_98[21:0];
  _RAND_99 = {1{`RANDOM}};
  _T_2207 = _RAND_99[21:0];
  _RAND_100 = {1{`RANDOM}};
  _T_2146 = _RAND_100[21:0];
  _RAND_101 = {1{`RANDOM}};
  _T_2085 = _RAND_101[21:0];
  _RAND_102 = {1{`RANDOM}};
  _T_2024 = _RAND_102[21:0];
  _RAND_103 = {1{`RANDOM}};
  _T_1963 = _RAND_103[21:0];
  _RAND_104 = {1{`RANDOM}};
  _T_1902 = _RAND_104[21:0];
  _RAND_105 = {1{`RANDOM}};
  _T_1841 = _RAND_105[21:0];
  _RAND_106 = {1{`RANDOM}};
  _T_1780 = _RAND_106[21:0];
  _RAND_107 = {1{`RANDOM}};
  _T_1719 = _RAND_107[21:0];
  _RAND_108 = {1{`RANDOM}};
  _T_1658 = _RAND_108[21:0];
  _RAND_109 = {1{`RANDOM}};
  _T_1597 = _RAND_109[21:0];
  _RAND_110 = {1{`RANDOM}};
  _T_1536 = _RAND_110[21:0];
  _RAND_111 = {1{`RANDOM}};
  _T_1475 = _RAND_111[21:0];
  _RAND_112 = {1{`RANDOM}};
  _T_1414 = _RAND_112[21:0];
  _RAND_113 = {1{`RANDOM}};
  _T_1353 = _RAND_113[21:0];
  _RAND_114 = {1{`RANDOM}};
  _T_1292 = _RAND_114[21:0];
  _RAND_115 = {1{`RANDOM}};
  _T_1231 = _RAND_115[21:0];
  _RAND_116 = {1{`RANDOM}};
  _T_1170 = _RAND_116[21:0];
  _RAND_117 = {1{`RANDOM}};
  _T_1109 = _RAND_117[21:0];
  _RAND_118 = {1{`RANDOM}};
  _T_1048 = _RAND_118[21:0];
  _RAND_119 = {1{`RANDOM}};
  _T_987 = _RAND_119[21:0];
  _RAND_120 = {1{`RANDOM}};
  _T_926 = _RAND_120[21:0];
  _RAND_121 = {1{`RANDOM}};
  _T_865 = _RAND_121[21:0];
  _RAND_122 = {1{`RANDOM}};
  _T_804 = _RAND_122[21:0];
  _RAND_123 = {1{`RANDOM}};
  _T_743 = _RAND_123[21:0];
  _RAND_124 = {1{`RANDOM}};
  _T_682 = _RAND_124[21:0];
  _RAND_125 = {1{`RANDOM}};
  _T_621 = _RAND_125[21:0];
  _RAND_126 = {1{`RANDOM}};
  _T_560 = _RAND_126[21:0];
  _RAND_127 = {1{`RANDOM}};
  _T_499 = _RAND_127[21:0];
  _RAND_128 = {1{`RANDOM}};
  _T_438 = _RAND_128[21:0];
  _RAND_129 = {1{`RANDOM}};
  _T_4303 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  _T_4242 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  _T_4181 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  _T_4120 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  _T_4059 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  _T_3998 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  _T_3937 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  _T_3876 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  _T_3815 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  _T_3754 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  _T_3693 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  _T_3632 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  _T_3571 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  _T_3510 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  _T_3449 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  _T_3388 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  _T_3327 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  _T_3266 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  _T_3205 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  _T_3144 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  _T_3083 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  _T_3022 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  _T_2961 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  _T_2900 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  _T_2839 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  _T_2778 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  _T_2717 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  _T_2656 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  _T_2595 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  _T_2534 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  _T_2473 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  _T_2412 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  _T_2351 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  _T_2290 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  _T_2229 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  _T_2168 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  _T_2107 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  _T_2046 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  _T_1985 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  _T_1924 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  _T_1863 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  _T_1802 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  _T_1741 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  _T_1680 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  _T_1619 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  _T_1558 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  _T_1497 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  _T_1436 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  _T_1375 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  _T_1314 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  _T_1253 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  _T_1192 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  _T_1131 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  _T_1070 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  _T_1009 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  _T_948 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  _T_887 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  _T_826 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  _T_765 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  _T_704 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  _T_643 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  _T_582 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  _T_521 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  _T_460 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  _T_4295 = _RAND_193[21:0];
  _RAND_194 = {1{`RANDOM}};
  _T_4234 = _RAND_194[21:0];
  _RAND_195 = {1{`RANDOM}};
  _T_4173 = _RAND_195[21:0];
  _RAND_196 = {1{`RANDOM}};
  _T_4112 = _RAND_196[21:0];
  _RAND_197 = {1{`RANDOM}};
  _T_4051 = _RAND_197[21:0];
  _RAND_198 = {1{`RANDOM}};
  _T_3990 = _RAND_198[21:0];
  _RAND_199 = {1{`RANDOM}};
  _T_3929 = _RAND_199[21:0];
  _RAND_200 = {1{`RANDOM}};
  _T_3868 = _RAND_200[21:0];
  _RAND_201 = {1{`RANDOM}};
  _T_3807 = _RAND_201[21:0];
  _RAND_202 = {1{`RANDOM}};
  _T_3746 = _RAND_202[21:0];
  _RAND_203 = {1{`RANDOM}};
  _T_3685 = _RAND_203[21:0];
  _RAND_204 = {1{`RANDOM}};
  _T_3624 = _RAND_204[21:0];
  _RAND_205 = {1{`RANDOM}};
  _T_3563 = _RAND_205[21:0];
  _RAND_206 = {1{`RANDOM}};
  _T_3502 = _RAND_206[21:0];
  _RAND_207 = {1{`RANDOM}};
  _T_3441 = _RAND_207[21:0];
  _RAND_208 = {1{`RANDOM}};
  _T_3380 = _RAND_208[21:0];
  _RAND_209 = {1{`RANDOM}};
  _T_3319 = _RAND_209[21:0];
  _RAND_210 = {1{`RANDOM}};
  _T_3258 = _RAND_210[21:0];
  _RAND_211 = {1{`RANDOM}};
  _T_3197 = _RAND_211[21:0];
  _RAND_212 = {1{`RANDOM}};
  _T_3136 = _RAND_212[21:0];
  _RAND_213 = {1{`RANDOM}};
  _T_3075 = _RAND_213[21:0];
  _RAND_214 = {1{`RANDOM}};
  _T_3014 = _RAND_214[21:0];
  _RAND_215 = {1{`RANDOM}};
  _T_2953 = _RAND_215[21:0];
  _RAND_216 = {1{`RANDOM}};
  _T_2892 = _RAND_216[21:0];
  _RAND_217 = {1{`RANDOM}};
  _T_2831 = _RAND_217[21:0];
  _RAND_218 = {1{`RANDOM}};
  _T_2770 = _RAND_218[21:0];
  _RAND_219 = {1{`RANDOM}};
  _T_2709 = _RAND_219[21:0];
  _RAND_220 = {1{`RANDOM}};
  _T_2648 = _RAND_220[21:0];
  _RAND_221 = {1{`RANDOM}};
  _T_2587 = _RAND_221[21:0];
  _RAND_222 = {1{`RANDOM}};
  _T_2526 = _RAND_222[21:0];
  _RAND_223 = {1{`RANDOM}};
  _T_2465 = _RAND_223[21:0];
  _RAND_224 = {1{`RANDOM}};
  _T_2404 = _RAND_224[21:0];
  _RAND_225 = {1{`RANDOM}};
  _T_2343 = _RAND_225[21:0];
  _RAND_226 = {1{`RANDOM}};
  _T_2282 = _RAND_226[21:0];
  _RAND_227 = {1{`RANDOM}};
  _T_2221 = _RAND_227[21:0];
  _RAND_228 = {1{`RANDOM}};
  _T_2160 = _RAND_228[21:0];
  _RAND_229 = {1{`RANDOM}};
  _T_2099 = _RAND_229[21:0];
  _RAND_230 = {1{`RANDOM}};
  _T_2038 = _RAND_230[21:0];
  _RAND_231 = {1{`RANDOM}};
  _T_1977 = _RAND_231[21:0];
  _RAND_232 = {1{`RANDOM}};
  _T_1916 = _RAND_232[21:0];
  _RAND_233 = {1{`RANDOM}};
  _T_1855 = _RAND_233[21:0];
  _RAND_234 = {1{`RANDOM}};
  _T_1794 = _RAND_234[21:0];
  _RAND_235 = {1{`RANDOM}};
  _T_1733 = _RAND_235[21:0];
  _RAND_236 = {1{`RANDOM}};
  _T_1672 = _RAND_236[21:0];
  _RAND_237 = {1{`RANDOM}};
  _T_1611 = _RAND_237[21:0];
  _RAND_238 = {1{`RANDOM}};
  _T_1550 = _RAND_238[21:0];
  _RAND_239 = {1{`RANDOM}};
  _T_1489 = _RAND_239[21:0];
  _RAND_240 = {1{`RANDOM}};
  _T_1428 = _RAND_240[21:0];
  _RAND_241 = {1{`RANDOM}};
  _T_1367 = _RAND_241[21:0];
  _RAND_242 = {1{`RANDOM}};
  _T_1306 = _RAND_242[21:0];
  _RAND_243 = {1{`RANDOM}};
  _T_1245 = _RAND_243[21:0];
  _RAND_244 = {1{`RANDOM}};
  _T_1184 = _RAND_244[21:0];
  _RAND_245 = {1{`RANDOM}};
  _T_1123 = _RAND_245[21:0];
  _RAND_246 = {1{`RANDOM}};
  _T_1062 = _RAND_246[21:0];
  _RAND_247 = {1{`RANDOM}};
  _T_1001 = _RAND_247[21:0];
  _RAND_248 = {1{`RANDOM}};
  _T_940 = _RAND_248[21:0];
  _RAND_249 = {1{`RANDOM}};
  _T_879 = _RAND_249[21:0];
  _RAND_250 = {1{`RANDOM}};
  _T_818 = _RAND_250[21:0];
  _RAND_251 = {1{`RANDOM}};
  _T_757 = _RAND_251[21:0];
  _RAND_252 = {1{`RANDOM}};
  _T_696 = _RAND_252[21:0];
  _RAND_253 = {1{`RANDOM}};
  _T_635 = _RAND_253[21:0];
  _RAND_254 = {1{`RANDOM}};
  _T_574 = _RAND_254[21:0];
  _RAND_255 = {1{`RANDOM}};
  _T_513 = _RAND_255[21:0];
  _RAND_256 = {1{`RANDOM}};
  _T_452 = _RAND_256[21:0];
  _RAND_257 = {1{`RANDOM}};
  _T_4317 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  _T_4256 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  _T_4195 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  _T_4134 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  _T_4073 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  _T_4012 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  _T_3951 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  _T_3890 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  _T_3829 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  _T_3768 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  _T_3707 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  _T_3646 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  _T_3585 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  _T_3524 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  _T_3463 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  _T_3402 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  _T_3341 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  _T_3280 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  _T_3219 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  _T_3158 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  _T_3097 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  _T_3036 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  _T_2975 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  _T_2914 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  _T_2853 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  _T_2792 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  _T_2731 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  _T_2670 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  _T_2609 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  _T_2548 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  _T_2487 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  _T_2426 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  _T_2365 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  _T_2304 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  _T_2243 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  _T_2182 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  _T_2121 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  _T_2060 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  _T_1999 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  _T_1938 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  _T_1877 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  _T_1816 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  _T_1755 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  _T_1694 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  _T_1633 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  _T_1572 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  _T_1511 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  _T_1450 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  _T_1389 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  _T_1328 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  _T_1267 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  _T_1206 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  _T_1145 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  _T_1084 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  _T_1023 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  _T_962 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  _T_901 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  _T_840 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  _T_779 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  _T_718 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  _T_657 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  _T_596 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  _T_535 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  _T_474 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  _T_4309 = _RAND_321[21:0];
  _RAND_322 = {1{`RANDOM}};
  _T_4248 = _RAND_322[21:0];
  _RAND_323 = {1{`RANDOM}};
  _T_4187 = _RAND_323[21:0];
  _RAND_324 = {1{`RANDOM}};
  _T_4126 = _RAND_324[21:0];
  _RAND_325 = {1{`RANDOM}};
  _T_4065 = _RAND_325[21:0];
  _RAND_326 = {1{`RANDOM}};
  _T_4004 = _RAND_326[21:0];
  _RAND_327 = {1{`RANDOM}};
  _T_3943 = _RAND_327[21:0];
  _RAND_328 = {1{`RANDOM}};
  _T_3882 = _RAND_328[21:0];
  _RAND_329 = {1{`RANDOM}};
  _T_3821 = _RAND_329[21:0];
  _RAND_330 = {1{`RANDOM}};
  _T_3760 = _RAND_330[21:0];
  _RAND_331 = {1{`RANDOM}};
  _T_3699 = _RAND_331[21:0];
  _RAND_332 = {1{`RANDOM}};
  _T_3638 = _RAND_332[21:0];
  _RAND_333 = {1{`RANDOM}};
  _T_3577 = _RAND_333[21:0];
  _RAND_334 = {1{`RANDOM}};
  _T_3516 = _RAND_334[21:0];
  _RAND_335 = {1{`RANDOM}};
  _T_3455 = _RAND_335[21:0];
  _RAND_336 = {1{`RANDOM}};
  _T_3394 = _RAND_336[21:0];
  _RAND_337 = {1{`RANDOM}};
  _T_3333 = _RAND_337[21:0];
  _RAND_338 = {1{`RANDOM}};
  _T_3272 = _RAND_338[21:0];
  _RAND_339 = {1{`RANDOM}};
  _T_3211 = _RAND_339[21:0];
  _RAND_340 = {1{`RANDOM}};
  _T_3150 = _RAND_340[21:0];
  _RAND_341 = {1{`RANDOM}};
  _T_3089 = _RAND_341[21:0];
  _RAND_342 = {1{`RANDOM}};
  _T_3028 = _RAND_342[21:0];
  _RAND_343 = {1{`RANDOM}};
  _T_2967 = _RAND_343[21:0];
  _RAND_344 = {1{`RANDOM}};
  _T_2906 = _RAND_344[21:0];
  _RAND_345 = {1{`RANDOM}};
  _T_2845 = _RAND_345[21:0];
  _RAND_346 = {1{`RANDOM}};
  _T_2784 = _RAND_346[21:0];
  _RAND_347 = {1{`RANDOM}};
  _T_2723 = _RAND_347[21:0];
  _RAND_348 = {1{`RANDOM}};
  _T_2662 = _RAND_348[21:0];
  _RAND_349 = {1{`RANDOM}};
  _T_2601 = _RAND_349[21:0];
  _RAND_350 = {1{`RANDOM}};
  _T_2540 = _RAND_350[21:0];
  _RAND_351 = {1{`RANDOM}};
  _T_2479 = _RAND_351[21:0];
  _RAND_352 = {1{`RANDOM}};
  _T_2418 = _RAND_352[21:0];
  _RAND_353 = {1{`RANDOM}};
  _T_2357 = _RAND_353[21:0];
  _RAND_354 = {1{`RANDOM}};
  _T_2296 = _RAND_354[21:0];
  _RAND_355 = {1{`RANDOM}};
  _T_2235 = _RAND_355[21:0];
  _RAND_356 = {1{`RANDOM}};
  _T_2174 = _RAND_356[21:0];
  _RAND_357 = {1{`RANDOM}};
  _T_2113 = _RAND_357[21:0];
  _RAND_358 = {1{`RANDOM}};
  _T_2052 = _RAND_358[21:0];
  _RAND_359 = {1{`RANDOM}};
  _T_1991 = _RAND_359[21:0];
  _RAND_360 = {1{`RANDOM}};
  _T_1930 = _RAND_360[21:0];
  _RAND_361 = {1{`RANDOM}};
  _T_1869 = _RAND_361[21:0];
  _RAND_362 = {1{`RANDOM}};
  _T_1808 = _RAND_362[21:0];
  _RAND_363 = {1{`RANDOM}};
  _T_1747 = _RAND_363[21:0];
  _RAND_364 = {1{`RANDOM}};
  _T_1686 = _RAND_364[21:0];
  _RAND_365 = {1{`RANDOM}};
  _T_1625 = _RAND_365[21:0];
  _RAND_366 = {1{`RANDOM}};
  _T_1564 = _RAND_366[21:0];
  _RAND_367 = {1{`RANDOM}};
  _T_1503 = _RAND_367[21:0];
  _RAND_368 = {1{`RANDOM}};
  _T_1442 = _RAND_368[21:0];
  _RAND_369 = {1{`RANDOM}};
  _T_1381 = _RAND_369[21:0];
  _RAND_370 = {1{`RANDOM}};
  _T_1320 = _RAND_370[21:0];
  _RAND_371 = {1{`RANDOM}};
  _T_1259 = _RAND_371[21:0];
  _RAND_372 = {1{`RANDOM}};
  _T_1198 = _RAND_372[21:0];
  _RAND_373 = {1{`RANDOM}};
  _T_1137 = _RAND_373[21:0];
  _RAND_374 = {1{`RANDOM}};
  _T_1076 = _RAND_374[21:0];
  _RAND_375 = {1{`RANDOM}};
  _T_1015 = _RAND_375[21:0];
  _RAND_376 = {1{`RANDOM}};
  _T_954 = _RAND_376[21:0];
  _RAND_377 = {1{`RANDOM}};
  _T_893 = _RAND_377[21:0];
  _RAND_378 = {1{`RANDOM}};
  _T_832 = _RAND_378[21:0];
  _RAND_379 = {1{`RANDOM}};
  _T_771 = _RAND_379[21:0];
  _RAND_380 = {1{`RANDOM}};
  _T_710 = _RAND_380[21:0];
  _RAND_381 = {1{`RANDOM}};
  _T_649 = _RAND_381[21:0];
  _RAND_382 = {1{`RANDOM}};
  _T_588 = _RAND_382[21:0];
  _RAND_383 = {1{`RANDOM}};
  _T_527 = _RAND_383[21:0];
  _RAND_384 = {1{`RANDOM}};
  _T_466 = _RAND_384[21:0];
  _RAND_385 = {1{`RANDOM}};
  _T_4331 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  _T_4270 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  _T_4209 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  _T_4148 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  _T_4087 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  _T_4026 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  _T_3965 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  _T_3904 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  _T_3843 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  _T_3782 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  _T_3721 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  _T_3660 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  _T_3599 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  _T_3538 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  _T_3477 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  _T_3416 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  _T_3355 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  _T_3294 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  _T_3233 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  _T_3172 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  _T_3111 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  _T_3050 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  _T_2989 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  _T_2928 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  _T_2867 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  _T_2806 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  _T_2745 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  _T_2684 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  _T_2623 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  _T_2562 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  _T_2501 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  _T_2440 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  _T_2379 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  _T_2318 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  _T_2257 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  _T_2196 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  _T_2135 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  _T_2074 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  _T_2013 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  _T_1952 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  _T_1891 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  _T_1830 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  _T_1769 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  _T_1708 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  _T_1647 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  _T_1586 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  _T_1525 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  _T_1464 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  _T_1403 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  _T_1342 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  _T_1281 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  _T_1220 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  _T_1159 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  _T_1098 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  _T_1037 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  _T_976 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  _T_915 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  _T_854 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  _T_793 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  _T_732 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  _T_671 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  _T_610 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  _T_549 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  _T_488 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  _T_4323 = _RAND_449[21:0];
  _RAND_450 = {1{`RANDOM}};
  _T_4262 = _RAND_450[21:0];
  _RAND_451 = {1{`RANDOM}};
  _T_4201 = _RAND_451[21:0];
  _RAND_452 = {1{`RANDOM}};
  _T_4140 = _RAND_452[21:0];
  _RAND_453 = {1{`RANDOM}};
  _T_4079 = _RAND_453[21:0];
  _RAND_454 = {1{`RANDOM}};
  _T_4018 = _RAND_454[21:0];
  _RAND_455 = {1{`RANDOM}};
  _T_3957 = _RAND_455[21:0];
  _RAND_456 = {1{`RANDOM}};
  _T_3896 = _RAND_456[21:0];
  _RAND_457 = {1{`RANDOM}};
  _T_3835 = _RAND_457[21:0];
  _RAND_458 = {1{`RANDOM}};
  _T_3774 = _RAND_458[21:0];
  _RAND_459 = {1{`RANDOM}};
  _T_3713 = _RAND_459[21:0];
  _RAND_460 = {1{`RANDOM}};
  _T_3652 = _RAND_460[21:0];
  _RAND_461 = {1{`RANDOM}};
  _T_3591 = _RAND_461[21:0];
  _RAND_462 = {1{`RANDOM}};
  _T_3530 = _RAND_462[21:0];
  _RAND_463 = {1{`RANDOM}};
  _T_3469 = _RAND_463[21:0];
  _RAND_464 = {1{`RANDOM}};
  _T_3408 = _RAND_464[21:0];
  _RAND_465 = {1{`RANDOM}};
  _T_3347 = _RAND_465[21:0];
  _RAND_466 = {1{`RANDOM}};
  _T_3286 = _RAND_466[21:0];
  _RAND_467 = {1{`RANDOM}};
  _T_3225 = _RAND_467[21:0];
  _RAND_468 = {1{`RANDOM}};
  _T_3164 = _RAND_468[21:0];
  _RAND_469 = {1{`RANDOM}};
  _T_3103 = _RAND_469[21:0];
  _RAND_470 = {1{`RANDOM}};
  _T_3042 = _RAND_470[21:0];
  _RAND_471 = {1{`RANDOM}};
  _T_2981 = _RAND_471[21:0];
  _RAND_472 = {1{`RANDOM}};
  _T_2920 = _RAND_472[21:0];
  _RAND_473 = {1{`RANDOM}};
  _T_2859 = _RAND_473[21:0];
  _RAND_474 = {1{`RANDOM}};
  _T_2798 = _RAND_474[21:0];
  _RAND_475 = {1{`RANDOM}};
  _T_2737 = _RAND_475[21:0];
  _RAND_476 = {1{`RANDOM}};
  _T_2676 = _RAND_476[21:0];
  _RAND_477 = {1{`RANDOM}};
  _T_2615 = _RAND_477[21:0];
  _RAND_478 = {1{`RANDOM}};
  _T_2554 = _RAND_478[21:0];
  _RAND_479 = {1{`RANDOM}};
  _T_2493 = _RAND_479[21:0];
  _RAND_480 = {1{`RANDOM}};
  _T_2432 = _RAND_480[21:0];
  _RAND_481 = {1{`RANDOM}};
  _T_2371 = _RAND_481[21:0];
  _RAND_482 = {1{`RANDOM}};
  _T_2310 = _RAND_482[21:0];
  _RAND_483 = {1{`RANDOM}};
  _T_2249 = _RAND_483[21:0];
  _RAND_484 = {1{`RANDOM}};
  _T_2188 = _RAND_484[21:0];
  _RAND_485 = {1{`RANDOM}};
  _T_2127 = _RAND_485[21:0];
  _RAND_486 = {1{`RANDOM}};
  _T_2066 = _RAND_486[21:0];
  _RAND_487 = {1{`RANDOM}};
  _T_2005 = _RAND_487[21:0];
  _RAND_488 = {1{`RANDOM}};
  _T_1944 = _RAND_488[21:0];
  _RAND_489 = {1{`RANDOM}};
  _T_1883 = _RAND_489[21:0];
  _RAND_490 = {1{`RANDOM}};
  _T_1822 = _RAND_490[21:0];
  _RAND_491 = {1{`RANDOM}};
  _T_1761 = _RAND_491[21:0];
  _RAND_492 = {1{`RANDOM}};
  _T_1700 = _RAND_492[21:0];
  _RAND_493 = {1{`RANDOM}};
  _T_1639 = _RAND_493[21:0];
  _RAND_494 = {1{`RANDOM}};
  _T_1578 = _RAND_494[21:0];
  _RAND_495 = {1{`RANDOM}};
  _T_1517 = _RAND_495[21:0];
  _RAND_496 = {1{`RANDOM}};
  _T_1456 = _RAND_496[21:0];
  _RAND_497 = {1{`RANDOM}};
  _T_1395 = _RAND_497[21:0];
  _RAND_498 = {1{`RANDOM}};
  _T_1334 = _RAND_498[21:0];
  _RAND_499 = {1{`RANDOM}};
  _T_1273 = _RAND_499[21:0];
  _RAND_500 = {1{`RANDOM}};
  _T_1212 = _RAND_500[21:0];
  _RAND_501 = {1{`RANDOM}};
  _T_1151 = _RAND_501[21:0];
  _RAND_502 = {1{`RANDOM}};
  _T_1090 = _RAND_502[21:0];
  _RAND_503 = {1{`RANDOM}};
  _T_1029 = _RAND_503[21:0];
  _RAND_504 = {1{`RANDOM}};
  _T_968 = _RAND_504[21:0];
  _RAND_505 = {1{`RANDOM}};
  _T_907 = _RAND_505[21:0];
  _RAND_506 = {1{`RANDOM}};
  _T_846 = _RAND_506[21:0];
  _RAND_507 = {1{`RANDOM}};
  _T_785 = _RAND_507[21:0];
  _RAND_508 = {1{`RANDOM}};
  _T_724 = _RAND_508[21:0];
  _RAND_509 = {1{`RANDOM}};
  _T_663 = _RAND_509[21:0];
  _RAND_510 = {1{`RANDOM}};
  _T_602 = _RAND_510[21:0];
  _RAND_511 = {1{`RANDOM}};
  _T_541 = _RAND_511[21:0];
  _RAND_512 = {1{`RANDOM}};
  _T_480 = _RAND_512[21:0];
  _RAND_513 = {1{`RANDOM}};
  _T_493 = _RAND_513[1:0];
  _RAND_514 = {1{`RANDOM}};
  _T_432 = _RAND_514[1:0];
  _RAND_515 = {1{`RANDOM}};
  _T_554 = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  _T_615 = _RAND_516[1:0];
  _RAND_517 = {1{`RANDOM}};
  _T_676 = _RAND_517[1:0];
  _RAND_518 = {1{`RANDOM}};
  _T_737 = _RAND_518[1:0];
  _RAND_519 = {1{`RANDOM}};
  _T_798 = _RAND_519[1:0];
  _RAND_520 = {1{`RANDOM}};
  _T_859 = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  _T_920 = _RAND_521[1:0];
  _RAND_522 = {1{`RANDOM}};
  _T_981 = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  _T_1042 = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  _T_1103 = _RAND_524[1:0];
  _RAND_525 = {1{`RANDOM}};
  _T_1164 = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  _T_1225 = _RAND_526[1:0];
  _RAND_527 = {1{`RANDOM}};
  _T_1286 = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  _T_1347 = _RAND_528[1:0];
  _RAND_529 = {1{`RANDOM}};
  _T_1408 = _RAND_529[1:0];
  _RAND_530 = {1{`RANDOM}};
  _T_1469 = _RAND_530[1:0];
  _RAND_531 = {1{`RANDOM}};
  _T_1530 = _RAND_531[1:0];
  _RAND_532 = {1{`RANDOM}};
  _T_1591 = _RAND_532[1:0];
  _RAND_533 = {1{`RANDOM}};
  _T_1652 = _RAND_533[1:0];
  _RAND_534 = {1{`RANDOM}};
  _T_1713 = _RAND_534[1:0];
  _RAND_535 = {1{`RANDOM}};
  _T_1774 = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  _T_1835 = _RAND_536[1:0];
  _RAND_537 = {1{`RANDOM}};
  _T_1896 = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  _T_1957 = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  _T_2018 = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  _T_2079 = _RAND_540[1:0];
  _RAND_541 = {1{`RANDOM}};
  _T_2140 = _RAND_541[1:0];
  _RAND_542 = {1{`RANDOM}};
  _T_2201 = _RAND_542[1:0];
  _RAND_543 = {1{`RANDOM}};
  _T_2262 = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  _T_2323 = _RAND_544[1:0];
  _RAND_545 = {1{`RANDOM}};
  _T_2384 = _RAND_545[1:0];
  _RAND_546 = {1{`RANDOM}};
  _T_2445 = _RAND_546[1:0];
  _RAND_547 = {1{`RANDOM}};
  _T_2506 = _RAND_547[1:0];
  _RAND_548 = {1{`RANDOM}};
  _T_2567 = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  _T_2628 = _RAND_549[1:0];
  _RAND_550 = {1{`RANDOM}};
  _T_2689 = _RAND_550[1:0];
  _RAND_551 = {1{`RANDOM}};
  _T_2750 = _RAND_551[1:0];
  _RAND_552 = {1{`RANDOM}};
  _T_2811 = _RAND_552[1:0];
  _RAND_553 = {1{`RANDOM}};
  _T_2872 = _RAND_553[1:0];
  _RAND_554 = {1{`RANDOM}};
  _T_2933 = _RAND_554[1:0];
  _RAND_555 = {1{`RANDOM}};
  _T_2994 = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  _T_3055 = _RAND_556[1:0];
  _RAND_557 = {1{`RANDOM}};
  _T_3116 = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  _T_3177 = _RAND_558[1:0];
  _RAND_559 = {1{`RANDOM}};
  _T_3238 = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  _T_3299 = _RAND_560[1:0];
  _RAND_561 = {1{`RANDOM}};
  _T_3360 = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  _T_3421 = _RAND_562[1:0];
  _RAND_563 = {1{`RANDOM}};
  _T_3482 = _RAND_563[1:0];
  _RAND_564 = {1{`RANDOM}};
  _T_3543 = _RAND_564[1:0];
  _RAND_565 = {1{`RANDOM}};
  _T_3604 = _RAND_565[1:0];
  _RAND_566 = {1{`RANDOM}};
  _T_3665 = _RAND_566[1:0];
  _RAND_567 = {1{`RANDOM}};
  _T_3726 = _RAND_567[1:0];
  _RAND_568 = {1{`RANDOM}};
  _T_3787 = _RAND_568[1:0];
  _RAND_569 = {1{`RANDOM}};
  _T_3848 = _RAND_569[1:0];
  _RAND_570 = {1{`RANDOM}};
  _T_3909 = _RAND_570[1:0];
  _RAND_571 = {1{`RANDOM}};
  _T_3970 = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  _T_4031 = _RAND_572[1:0];
  _RAND_573 = {1{`RANDOM}};
  _T_4092 = _RAND_573[1:0];
  _RAND_574 = {1{`RANDOM}};
  _T_4153 = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  _T_4214 = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  _T_4275 = _RAND_576[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_4 <= 2'h0;
    end else if (_T_15) begin
      if (io_block) begin
        _T_4 <= 2'h3;
      end else begin
        _T_4 <= 2'h0;
      end
    end else if (_T_13) begin
      if (io_block) begin
        _T_4 <= 2'h3;
      end else begin
        _T_4 <= 2'h0;
      end
    end else if (_T_11) begin
      if (io_cacheOut_r_last_i) begin
        _T_4 <= 2'h0;
      end else begin
        _T_4 <= 2'h1;
      end
    end else if (io_cacheIn_valid) begin
      if (_T_286) begin
        _T_4 <= 2'h2;
      end else begin
        _T_4 <= 2'h1;
      end
    end else begin
      _T_4 <= 2'h0;
    end
    if (_T_440) begin
      _T_4289 <= 1'h0;
    end else begin
      _T_4289 <= _GEN_569;
    end
    if (_T_440) begin
      _T_4228 <= 1'h0;
    end else begin
      _T_4228 <= _GEN_560;
    end
    if (_T_440) begin
      _T_4167 <= 1'h0;
    end else begin
      _T_4167 <= _GEN_551;
    end
    if (_T_440) begin
      _T_4106 <= 1'h0;
    end else begin
      _T_4106 <= _GEN_542;
    end
    if (_T_440) begin
      _T_4045 <= 1'h0;
    end else begin
      _T_4045 <= _GEN_533;
    end
    if (_T_440) begin
      _T_3984 <= 1'h0;
    end else begin
      _T_3984 <= _GEN_524;
    end
    if (_T_440) begin
      _T_3923 <= 1'h0;
    end else begin
      _T_3923 <= _GEN_515;
    end
    if (_T_440) begin
      _T_3862 <= 1'h0;
    end else begin
      _T_3862 <= _GEN_506;
    end
    if (_T_440) begin
      _T_3801 <= 1'h0;
    end else begin
      _T_3801 <= _GEN_497;
    end
    if (_T_440) begin
      _T_3740 <= 1'h0;
    end else begin
      _T_3740 <= _GEN_488;
    end
    if (_T_440) begin
      _T_3679 <= 1'h0;
    end else begin
      _T_3679 <= _GEN_479;
    end
    if (_T_440) begin
      _T_3618 <= 1'h0;
    end else begin
      _T_3618 <= _GEN_470;
    end
    if (_T_440) begin
      _T_3557 <= 1'h0;
    end else begin
      _T_3557 <= _GEN_461;
    end
    if (_T_440) begin
      _T_3496 <= 1'h0;
    end else begin
      _T_3496 <= _GEN_452;
    end
    if (_T_440) begin
      _T_3435 <= 1'h0;
    end else begin
      _T_3435 <= _GEN_443;
    end
    if (_T_440) begin
      _T_3374 <= 1'h0;
    end else begin
      _T_3374 <= _GEN_434;
    end
    if (_T_440) begin
      _T_3313 <= 1'h0;
    end else begin
      _T_3313 <= _GEN_425;
    end
    if (_T_440) begin
      _T_3252 <= 1'h0;
    end else begin
      _T_3252 <= _GEN_416;
    end
    if (_T_440) begin
      _T_3191 <= 1'h0;
    end else begin
      _T_3191 <= _GEN_407;
    end
    if (_T_440) begin
      _T_3130 <= 1'h0;
    end else begin
      _T_3130 <= _GEN_398;
    end
    if (_T_440) begin
      _T_3069 <= 1'h0;
    end else begin
      _T_3069 <= _GEN_389;
    end
    if (_T_440) begin
      _T_3008 <= 1'h0;
    end else begin
      _T_3008 <= _GEN_380;
    end
    if (_T_440) begin
      _T_2947 <= 1'h0;
    end else begin
      _T_2947 <= _GEN_371;
    end
    if (_T_440) begin
      _T_2886 <= 1'h0;
    end else begin
      _T_2886 <= _GEN_362;
    end
    if (_T_440) begin
      _T_2825 <= 1'h0;
    end else begin
      _T_2825 <= _GEN_353;
    end
    if (_T_440) begin
      _T_2764 <= 1'h0;
    end else begin
      _T_2764 <= _GEN_344;
    end
    if (_T_440) begin
      _T_2703 <= 1'h0;
    end else begin
      _T_2703 <= _GEN_335;
    end
    if (_T_440) begin
      _T_2642 <= 1'h0;
    end else begin
      _T_2642 <= _GEN_326;
    end
    if (_T_440) begin
      _T_2581 <= 1'h0;
    end else begin
      _T_2581 <= _GEN_317;
    end
    if (_T_440) begin
      _T_2520 <= 1'h0;
    end else begin
      _T_2520 <= _GEN_308;
    end
    if (_T_440) begin
      _T_2459 <= 1'h0;
    end else begin
      _T_2459 <= _GEN_299;
    end
    if (_T_440) begin
      _T_2398 <= 1'h0;
    end else begin
      _T_2398 <= _GEN_290;
    end
    if (_T_440) begin
      _T_2337 <= 1'h0;
    end else begin
      _T_2337 <= _GEN_281;
    end
    if (_T_440) begin
      _T_2276 <= 1'h0;
    end else begin
      _T_2276 <= _GEN_272;
    end
    if (_T_440) begin
      _T_2215 <= 1'h0;
    end else begin
      _T_2215 <= _GEN_263;
    end
    if (_T_440) begin
      _T_2154 <= 1'h0;
    end else begin
      _T_2154 <= _GEN_254;
    end
    if (_T_440) begin
      _T_2093 <= 1'h0;
    end else begin
      _T_2093 <= _GEN_245;
    end
    if (_T_440) begin
      _T_2032 <= 1'h0;
    end else begin
      _T_2032 <= _GEN_236;
    end
    if (_T_440) begin
      _T_1971 <= 1'h0;
    end else begin
      _T_1971 <= _GEN_227;
    end
    if (_T_440) begin
      _T_1910 <= 1'h0;
    end else begin
      _T_1910 <= _GEN_218;
    end
    if (_T_440) begin
      _T_1849 <= 1'h0;
    end else begin
      _T_1849 <= _GEN_209;
    end
    if (_T_440) begin
      _T_1788 <= 1'h0;
    end else begin
      _T_1788 <= _GEN_200;
    end
    if (_T_440) begin
      _T_1727 <= 1'h0;
    end else begin
      _T_1727 <= _GEN_191;
    end
    if (_T_440) begin
      _T_1666 <= 1'h0;
    end else begin
      _T_1666 <= _GEN_182;
    end
    if (_T_440) begin
      _T_1605 <= 1'h0;
    end else begin
      _T_1605 <= _GEN_173;
    end
    if (_T_440) begin
      _T_1544 <= 1'h0;
    end else begin
      _T_1544 <= _GEN_164;
    end
    if (_T_440) begin
      _T_1483 <= 1'h0;
    end else begin
      _T_1483 <= _GEN_155;
    end
    if (_T_440) begin
      _T_1422 <= 1'h0;
    end else begin
      _T_1422 <= _GEN_146;
    end
    if (_T_440) begin
      _T_1361 <= 1'h0;
    end else begin
      _T_1361 <= _GEN_137;
    end
    if (_T_440) begin
      _T_1300 <= 1'h0;
    end else begin
      _T_1300 <= _GEN_128;
    end
    if (_T_440) begin
      _T_1239 <= 1'h0;
    end else begin
      _T_1239 <= _GEN_119;
    end
    if (_T_440) begin
      _T_1178 <= 1'h0;
    end else begin
      _T_1178 <= _GEN_110;
    end
    if (_T_440) begin
      _T_1117 <= 1'h0;
    end else begin
      _T_1117 <= _GEN_101;
    end
    if (_T_440) begin
      _T_1056 <= 1'h0;
    end else begin
      _T_1056 <= _GEN_92;
    end
    if (_T_440) begin
      _T_995 <= 1'h0;
    end else begin
      _T_995 <= _GEN_83;
    end
    if (_T_440) begin
      _T_934 <= 1'h0;
    end else begin
      _T_934 <= _GEN_74;
    end
    if (_T_440) begin
      _T_873 <= 1'h0;
    end else begin
      _T_873 <= _GEN_65;
    end
    if (_T_440) begin
      _T_812 <= 1'h0;
    end else begin
      _T_812 <= _GEN_56;
    end
    if (_T_440) begin
      _T_751 <= 1'h0;
    end else begin
      _T_751 <= _GEN_47;
    end
    if (_T_440) begin
      _T_690 <= 1'h0;
    end else begin
      _T_690 <= _GEN_38;
    end
    if (_T_440) begin
      _T_629 <= 1'h0;
    end else begin
      _T_629 <= _GEN_29;
    end
    if (_T_440) begin
      _T_568 <= 1'h0;
    end else begin
      _T_568 <= _GEN_20;
    end
    if (_T_440) begin
      _T_507 <= 1'h0;
    end else begin
      _T_507 <= _GEN_11;
    end
    if (_T_440) begin
      _T_446 <= 1'h0;
    end else begin
      _T_446 <= _GEN_2;
    end
    if (reset) begin
      _T_4281 <= 22'h0;
    end else if (_T_4280) begin
      _T_4281 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4220 <= 22'h0;
    end else if (_T_4219) begin
      _T_4220 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4159 <= 22'h0;
    end else if (_T_4158) begin
      _T_4159 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4098 <= 22'h0;
    end else if (_T_4097) begin
      _T_4098 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4037 <= 22'h0;
    end else if (_T_4036) begin
      _T_4037 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3976 <= 22'h0;
    end else if (_T_3975) begin
      _T_3976 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3915 <= 22'h0;
    end else if (_T_3914) begin
      _T_3915 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3854 <= 22'h0;
    end else if (_T_3853) begin
      _T_3854 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3793 <= 22'h0;
    end else if (_T_3792) begin
      _T_3793 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3732 <= 22'h0;
    end else if (_T_3731) begin
      _T_3732 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3671 <= 22'h0;
    end else if (_T_3670) begin
      _T_3671 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3610 <= 22'h0;
    end else if (_T_3609) begin
      _T_3610 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3549 <= 22'h0;
    end else if (_T_3548) begin
      _T_3549 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3488 <= 22'h0;
    end else if (_T_3487) begin
      _T_3488 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3427 <= 22'h0;
    end else if (_T_3426) begin
      _T_3427 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3366 <= 22'h0;
    end else if (_T_3365) begin
      _T_3366 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3305 <= 22'h0;
    end else if (_T_3304) begin
      _T_3305 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3244 <= 22'h0;
    end else if (_T_3243) begin
      _T_3244 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3183 <= 22'h0;
    end else if (_T_3182) begin
      _T_3183 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3122 <= 22'h0;
    end else if (_T_3121) begin
      _T_3122 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3061 <= 22'h0;
    end else if (_T_3060) begin
      _T_3061 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3000 <= 22'h0;
    end else if (_T_2999) begin
      _T_3000 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2939 <= 22'h0;
    end else if (_T_2938) begin
      _T_2939 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2878 <= 22'h0;
    end else if (_T_2877) begin
      _T_2878 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2817 <= 22'h0;
    end else if (_T_2816) begin
      _T_2817 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2756 <= 22'h0;
    end else if (_T_2755) begin
      _T_2756 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2695 <= 22'h0;
    end else if (_T_2694) begin
      _T_2695 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2634 <= 22'h0;
    end else if (_T_2633) begin
      _T_2634 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2573 <= 22'h0;
    end else if (_T_2572) begin
      _T_2573 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2512 <= 22'h0;
    end else if (_T_2511) begin
      _T_2512 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2451 <= 22'h0;
    end else if (_T_2450) begin
      _T_2451 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2390 <= 22'h0;
    end else if (_T_2389) begin
      _T_2390 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2329 <= 22'h0;
    end else if (_T_2328) begin
      _T_2329 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2268 <= 22'h0;
    end else if (_T_2267) begin
      _T_2268 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2207 <= 22'h0;
    end else if (_T_2206) begin
      _T_2207 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2146 <= 22'h0;
    end else if (_T_2145) begin
      _T_2146 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2085 <= 22'h0;
    end else if (_T_2084) begin
      _T_2085 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2024 <= 22'h0;
    end else if (_T_2023) begin
      _T_2024 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1963 <= 22'h0;
    end else if (_T_1962) begin
      _T_1963 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1902 <= 22'h0;
    end else if (_T_1901) begin
      _T_1902 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1841 <= 22'h0;
    end else if (_T_1840) begin
      _T_1841 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1780 <= 22'h0;
    end else if (_T_1779) begin
      _T_1780 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1719 <= 22'h0;
    end else if (_T_1718) begin
      _T_1719 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1658 <= 22'h0;
    end else if (_T_1657) begin
      _T_1658 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1597 <= 22'h0;
    end else if (_T_1596) begin
      _T_1597 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1536 <= 22'h0;
    end else if (_T_1535) begin
      _T_1536 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1475 <= 22'h0;
    end else if (_T_1474) begin
      _T_1475 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1414 <= 22'h0;
    end else if (_T_1413) begin
      _T_1414 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1353 <= 22'h0;
    end else if (_T_1352) begin
      _T_1353 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1292 <= 22'h0;
    end else if (_T_1291) begin
      _T_1292 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1231 <= 22'h0;
    end else if (_T_1230) begin
      _T_1231 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1170 <= 22'h0;
    end else if (_T_1169) begin
      _T_1170 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1109 <= 22'h0;
    end else if (_T_1108) begin
      _T_1109 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1048 <= 22'h0;
    end else if (_T_1047) begin
      _T_1048 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_987 <= 22'h0;
    end else if (_T_986) begin
      _T_987 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_926 <= 22'h0;
    end else if (_T_925) begin
      _T_926 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_865 <= 22'h0;
    end else if (_T_864) begin
      _T_865 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_804 <= 22'h0;
    end else if (_T_803) begin
      _T_804 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_743 <= 22'h0;
    end else if (_T_742) begin
      _T_743 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_682 <= 22'h0;
    end else if (_T_681) begin
      _T_682 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_621 <= 22'h0;
    end else if (_T_620) begin
      _T_621 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_560 <= 22'h0;
    end else if (_T_559) begin
      _T_560 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_499 <= 22'h0;
    end else if (_T_498) begin
      _T_499 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_438 <= 22'h0;
    end else if (_T_437) begin
      _T_438 <= io_cacheIn_addr[31:10];
    end
    if (_T_440) begin
      _T_4303 <= 1'h0;
    end else begin
      _T_4303 <= _GEN_571;
    end
    if (_T_440) begin
      _T_4242 <= 1'h0;
    end else begin
      _T_4242 <= _GEN_562;
    end
    if (_T_440) begin
      _T_4181 <= 1'h0;
    end else begin
      _T_4181 <= _GEN_553;
    end
    if (_T_440) begin
      _T_4120 <= 1'h0;
    end else begin
      _T_4120 <= _GEN_544;
    end
    if (_T_440) begin
      _T_4059 <= 1'h0;
    end else begin
      _T_4059 <= _GEN_535;
    end
    if (_T_440) begin
      _T_3998 <= 1'h0;
    end else begin
      _T_3998 <= _GEN_526;
    end
    if (_T_440) begin
      _T_3937 <= 1'h0;
    end else begin
      _T_3937 <= _GEN_517;
    end
    if (_T_440) begin
      _T_3876 <= 1'h0;
    end else begin
      _T_3876 <= _GEN_508;
    end
    if (_T_440) begin
      _T_3815 <= 1'h0;
    end else begin
      _T_3815 <= _GEN_499;
    end
    if (_T_440) begin
      _T_3754 <= 1'h0;
    end else begin
      _T_3754 <= _GEN_490;
    end
    if (_T_440) begin
      _T_3693 <= 1'h0;
    end else begin
      _T_3693 <= _GEN_481;
    end
    if (_T_440) begin
      _T_3632 <= 1'h0;
    end else begin
      _T_3632 <= _GEN_472;
    end
    if (_T_440) begin
      _T_3571 <= 1'h0;
    end else begin
      _T_3571 <= _GEN_463;
    end
    if (_T_440) begin
      _T_3510 <= 1'h0;
    end else begin
      _T_3510 <= _GEN_454;
    end
    if (_T_440) begin
      _T_3449 <= 1'h0;
    end else begin
      _T_3449 <= _GEN_445;
    end
    if (_T_440) begin
      _T_3388 <= 1'h0;
    end else begin
      _T_3388 <= _GEN_436;
    end
    if (_T_440) begin
      _T_3327 <= 1'h0;
    end else begin
      _T_3327 <= _GEN_427;
    end
    if (_T_440) begin
      _T_3266 <= 1'h0;
    end else begin
      _T_3266 <= _GEN_418;
    end
    if (_T_440) begin
      _T_3205 <= 1'h0;
    end else begin
      _T_3205 <= _GEN_409;
    end
    if (_T_440) begin
      _T_3144 <= 1'h0;
    end else begin
      _T_3144 <= _GEN_400;
    end
    if (_T_440) begin
      _T_3083 <= 1'h0;
    end else begin
      _T_3083 <= _GEN_391;
    end
    if (_T_440) begin
      _T_3022 <= 1'h0;
    end else begin
      _T_3022 <= _GEN_382;
    end
    if (_T_440) begin
      _T_2961 <= 1'h0;
    end else begin
      _T_2961 <= _GEN_373;
    end
    if (_T_440) begin
      _T_2900 <= 1'h0;
    end else begin
      _T_2900 <= _GEN_364;
    end
    if (_T_440) begin
      _T_2839 <= 1'h0;
    end else begin
      _T_2839 <= _GEN_355;
    end
    if (_T_440) begin
      _T_2778 <= 1'h0;
    end else begin
      _T_2778 <= _GEN_346;
    end
    if (_T_440) begin
      _T_2717 <= 1'h0;
    end else begin
      _T_2717 <= _GEN_337;
    end
    if (_T_440) begin
      _T_2656 <= 1'h0;
    end else begin
      _T_2656 <= _GEN_328;
    end
    if (_T_440) begin
      _T_2595 <= 1'h0;
    end else begin
      _T_2595 <= _GEN_319;
    end
    if (_T_440) begin
      _T_2534 <= 1'h0;
    end else begin
      _T_2534 <= _GEN_310;
    end
    if (_T_440) begin
      _T_2473 <= 1'h0;
    end else begin
      _T_2473 <= _GEN_301;
    end
    if (_T_440) begin
      _T_2412 <= 1'h0;
    end else begin
      _T_2412 <= _GEN_292;
    end
    if (_T_440) begin
      _T_2351 <= 1'h0;
    end else begin
      _T_2351 <= _GEN_283;
    end
    if (_T_440) begin
      _T_2290 <= 1'h0;
    end else begin
      _T_2290 <= _GEN_274;
    end
    if (_T_440) begin
      _T_2229 <= 1'h0;
    end else begin
      _T_2229 <= _GEN_265;
    end
    if (_T_440) begin
      _T_2168 <= 1'h0;
    end else begin
      _T_2168 <= _GEN_256;
    end
    if (_T_440) begin
      _T_2107 <= 1'h0;
    end else begin
      _T_2107 <= _GEN_247;
    end
    if (_T_440) begin
      _T_2046 <= 1'h0;
    end else begin
      _T_2046 <= _GEN_238;
    end
    if (_T_440) begin
      _T_1985 <= 1'h0;
    end else begin
      _T_1985 <= _GEN_229;
    end
    if (_T_440) begin
      _T_1924 <= 1'h0;
    end else begin
      _T_1924 <= _GEN_220;
    end
    if (_T_440) begin
      _T_1863 <= 1'h0;
    end else begin
      _T_1863 <= _GEN_211;
    end
    if (_T_440) begin
      _T_1802 <= 1'h0;
    end else begin
      _T_1802 <= _GEN_202;
    end
    if (_T_440) begin
      _T_1741 <= 1'h0;
    end else begin
      _T_1741 <= _GEN_193;
    end
    if (_T_440) begin
      _T_1680 <= 1'h0;
    end else begin
      _T_1680 <= _GEN_184;
    end
    if (_T_440) begin
      _T_1619 <= 1'h0;
    end else begin
      _T_1619 <= _GEN_175;
    end
    if (_T_440) begin
      _T_1558 <= 1'h0;
    end else begin
      _T_1558 <= _GEN_166;
    end
    if (_T_440) begin
      _T_1497 <= 1'h0;
    end else begin
      _T_1497 <= _GEN_157;
    end
    if (_T_440) begin
      _T_1436 <= 1'h0;
    end else begin
      _T_1436 <= _GEN_148;
    end
    if (_T_440) begin
      _T_1375 <= 1'h0;
    end else begin
      _T_1375 <= _GEN_139;
    end
    if (_T_440) begin
      _T_1314 <= 1'h0;
    end else begin
      _T_1314 <= _GEN_130;
    end
    if (_T_440) begin
      _T_1253 <= 1'h0;
    end else begin
      _T_1253 <= _GEN_121;
    end
    if (_T_440) begin
      _T_1192 <= 1'h0;
    end else begin
      _T_1192 <= _GEN_112;
    end
    if (_T_440) begin
      _T_1131 <= 1'h0;
    end else begin
      _T_1131 <= _GEN_103;
    end
    if (_T_440) begin
      _T_1070 <= 1'h0;
    end else begin
      _T_1070 <= _GEN_94;
    end
    if (_T_440) begin
      _T_1009 <= 1'h0;
    end else begin
      _T_1009 <= _GEN_85;
    end
    if (_T_440) begin
      _T_948 <= 1'h0;
    end else begin
      _T_948 <= _GEN_76;
    end
    if (_T_440) begin
      _T_887 <= 1'h0;
    end else begin
      _T_887 <= _GEN_67;
    end
    if (_T_440) begin
      _T_826 <= 1'h0;
    end else begin
      _T_826 <= _GEN_58;
    end
    if (_T_440) begin
      _T_765 <= 1'h0;
    end else begin
      _T_765 <= _GEN_49;
    end
    if (_T_440) begin
      _T_704 <= 1'h0;
    end else begin
      _T_704 <= _GEN_40;
    end
    if (_T_440) begin
      _T_643 <= 1'h0;
    end else begin
      _T_643 <= _GEN_31;
    end
    if (_T_440) begin
      _T_582 <= 1'h0;
    end else begin
      _T_582 <= _GEN_22;
    end
    if (_T_440) begin
      _T_521 <= 1'h0;
    end else begin
      _T_521 <= _GEN_13;
    end
    if (_T_440) begin
      _T_460 <= 1'h0;
    end else begin
      _T_460 <= _GEN_4;
    end
    if (reset) begin
      _T_4295 <= 22'h0;
    end else if (_T_4294) begin
      _T_4295 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4234 <= 22'h0;
    end else if (_T_4233) begin
      _T_4234 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4173 <= 22'h0;
    end else if (_T_4172) begin
      _T_4173 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4112 <= 22'h0;
    end else if (_T_4111) begin
      _T_4112 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4051 <= 22'h0;
    end else if (_T_4050) begin
      _T_4051 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3990 <= 22'h0;
    end else if (_T_3989) begin
      _T_3990 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3929 <= 22'h0;
    end else if (_T_3928) begin
      _T_3929 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3868 <= 22'h0;
    end else if (_T_3867) begin
      _T_3868 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3807 <= 22'h0;
    end else if (_T_3806) begin
      _T_3807 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3746 <= 22'h0;
    end else if (_T_3745) begin
      _T_3746 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3685 <= 22'h0;
    end else if (_T_3684) begin
      _T_3685 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3624 <= 22'h0;
    end else if (_T_3623) begin
      _T_3624 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3563 <= 22'h0;
    end else if (_T_3562) begin
      _T_3563 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3502 <= 22'h0;
    end else if (_T_3501) begin
      _T_3502 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3441 <= 22'h0;
    end else if (_T_3440) begin
      _T_3441 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3380 <= 22'h0;
    end else if (_T_3379) begin
      _T_3380 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3319 <= 22'h0;
    end else if (_T_3318) begin
      _T_3319 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3258 <= 22'h0;
    end else if (_T_3257) begin
      _T_3258 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3197 <= 22'h0;
    end else if (_T_3196) begin
      _T_3197 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3136 <= 22'h0;
    end else if (_T_3135) begin
      _T_3136 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3075 <= 22'h0;
    end else if (_T_3074) begin
      _T_3075 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3014 <= 22'h0;
    end else if (_T_3013) begin
      _T_3014 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2953 <= 22'h0;
    end else if (_T_2952) begin
      _T_2953 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2892 <= 22'h0;
    end else if (_T_2891) begin
      _T_2892 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2831 <= 22'h0;
    end else if (_T_2830) begin
      _T_2831 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2770 <= 22'h0;
    end else if (_T_2769) begin
      _T_2770 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2709 <= 22'h0;
    end else if (_T_2708) begin
      _T_2709 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2648 <= 22'h0;
    end else if (_T_2647) begin
      _T_2648 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2587 <= 22'h0;
    end else if (_T_2586) begin
      _T_2587 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2526 <= 22'h0;
    end else if (_T_2525) begin
      _T_2526 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2465 <= 22'h0;
    end else if (_T_2464) begin
      _T_2465 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2404 <= 22'h0;
    end else if (_T_2403) begin
      _T_2404 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2343 <= 22'h0;
    end else if (_T_2342) begin
      _T_2343 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2282 <= 22'h0;
    end else if (_T_2281) begin
      _T_2282 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2221 <= 22'h0;
    end else if (_T_2220) begin
      _T_2221 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2160 <= 22'h0;
    end else if (_T_2159) begin
      _T_2160 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2099 <= 22'h0;
    end else if (_T_2098) begin
      _T_2099 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2038 <= 22'h0;
    end else if (_T_2037) begin
      _T_2038 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1977 <= 22'h0;
    end else if (_T_1976) begin
      _T_1977 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1916 <= 22'h0;
    end else if (_T_1915) begin
      _T_1916 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1855 <= 22'h0;
    end else if (_T_1854) begin
      _T_1855 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1794 <= 22'h0;
    end else if (_T_1793) begin
      _T_1794 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1733 <= 22'h0;
    end else if (_T_1732) begin
      _T_1733 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1672 <= 22'h0;
    end else if (_T_1671) begin
      _T_1672 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1611 <= 22'h0;
    end else if (_T_1610) begin
      _T_1611 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1550 <= 22'h0;
    end else if (_T_1549) begin
      _T_1550 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1489 <= 22'h0;
    end else if (_T_1488) begin
      _T_1489 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1428 <= 22'h0;
    end else if (_T_1427) begin
      _T_1428 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1367 <= 22'h0;
    end else if (_T_1366) begin
      _T_1367 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1306 <= 22'h0;
    end else if (_T_1305) begin
      _T_1306 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1245 <= 22'h0;
    end else if (_T_1244) begin
      _T_1245 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1184 <= 22'h0;
    end else if (_T_1183) begin
      _T_1184 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1123 <= 22'h0;
    end else if (_T_1122) begin
      _T_1123 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1062 <= 22'h0;
    end else if (_T_1061) begin
      _T_1062 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1001 <= 22'h0;
    end else if (_T_1000) begin
      _T_1001 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_940 <= 22'h0;
    end else if (_T_939) begin
      _T_940 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_879 <= 22'h0;
    end else if (_T_878) begin
      _T_879 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_818 <= 22'h0;
    end else if (_T_817) begin
      _T_818 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_757 <= 22'h0;
    end else if (_T_756) begin
      _T_757 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_696 <= 22'h0;
    end else if (_T_695) begin
      _T_696 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_635 <= 22'h0;
    end else if (_T_634) begin
      _T_635 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_574 <= 22'h0;
    end else if (_T_573) begin
      _T_574 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_513 <= 22'h0;
    end else if (_T_512) begin
      _T_513 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_452 <= 22'h0;
    end else if (_T_451) begin
      _T_452 <= io_cacheIn_addr[31:10];
    end
    if (_T_440) begin
      _T_4317 <= 1'h0;
    end else begin
      _T_4317 <= _GEN_573;
    end
    if (_T_440) begin
      _T_4256 <= 1'h0;
    end else begin
      _T_4256 <= _GEN_564;
    end
    if (_T_440) begin
      _T_4195 <= 1'h0;
    end else begin
      _T_4195 <= _GEN_555;
    end
    if (_T_440) begin
      _T_4134 <= 1'h0;
    end else begin
      _T_4134 <= _GEN_546;
    end
    if (_T_440) begin
      _T_4073 <= 1'h0;
    end else begin
      _T_4073 <= _GEN_537;
    end
    if (_T_440) begin
      _T_4012 <= 1'h0;
    end else begin
      _T_4012 <= _GEN_528;
    end
    if (_T_440) begin
      _T_3951 <= 1'h0;
    end else begin
      _T_3951 <= _GEN_519;
    end
    if (_T_440) begin
      _T_3890 <= 1'h0;
    end else begin
      _T_3890 <= _GEN_510;
    end
    if (_T_440) begin
      _T_3829 <= 1'h0;
    end else begin
      _T_3829 <= _GEN_501;
    end
    if (_T_440) begin
      _T_3768 <= 1'h0;
    end else begin
      _T_3768 <= _GEN_492;
    end
    if (_T_440) begin
      _T_3707 <= 1'h0;
    end else begin
      _T_3707 <= _GEN_483;
    end
    if (_T_440) begin
      _T_3646 <= 1'h0;
    end else begin
      _T_3646 <= _GEN_474;
    end
    if (_T_440) begin
      _T_3585 <= 1'h0;
    end else begin
      _T_3585 <= _GEN_465;
    end
    if (_T_440) begin
      _T_3524 <= 1'h0;
    end else begin
      _T_3524 <= _GEN_456;
    end
    if (_T_440) begin
      _T_3463 <= 1'h0;
    end else begin
      _T_3463 <= _GEN_447;
    end
    if (_T_440) begin
      _T_3402 <= 1'h0;
    end else begin
      _T_3402 <= _GEN_438;
    end
    if (_T_440) begin
      _T_3341 <= 1'h0;
    end else begin
      _T_3341 <= _GEN_429;
    end
    if (_T_440) begin
      _T_3280 <= 1'h0;
    end else begin
      _T_3280 <= _GEN_420;
    end
    if (_T_440) begin
      _T_3219 <= 1'h0;
    end else begin
      _T_3219 <= _GEN_411;
    end
    if (_T_440) begin
      _T_3158 <= 1'h0;
    end else begin
      _T_3158 <= _GEN_402;
    end
    if (_T_440) begin
      _T_3097 <= 1'h0;
    end else begin
      _T_3097 <= _GEN_393;
    end
    if (_T_440) begin
      _T_3036 <= 1'h0;
    end else begin
      _T_3036 <= _GEN_384;
    end
    if (_T_440) begin
      _T_2975 <= 1'h0;
    end else begin
      _T_2975 <= _GEN_375;
    end
    if (_T_440) begin
      _T_2914 <= 1'h0;
    end else begin
      _T_2914 <= _GEN_366;
    end
    if (_T_440) begin
      _T_2853 <= 1'h0;
    end else begin
      _T_2853 <= _GEN_357;
    end
    if (_T_440) begin
      _T_2792 <= 1'h0;
    end else begin
      _T_2792 <= _GEN_348;
    end
    if (_T_440) begin
      _T_2731 <= 1'h0;
    end else begin
      _T_2731 <= _GEN_339;
    end
    if (_T_440) begin
      _T_2670 <= 1'h0;
    end else begin
      _T_2670 <= _GEN_330;
    end
    if (_T_440) begin
      _T_2609 <= 1'h0;
    end else begin
      _T_2609 <= _GEN_321;
    end
    if (_T_440) begin
      _T_2548 <= 1'h0;
    end else begin
      _T_2548 <= _GEN_312;
    end
    if (_T_440) begin
      _T_2487 <= 1'h0;
    end else begin
      _T_2487 <= _GEN_303;
    end
    if (_T_440) begin
      _T_2426 <= 1'h0;
    end else begin
      _T_2426 <= _GEN_294;
    end
    if (_T_440) begin
      _T_2365 <= 1'h0;
    end else begin
      _T_2365 <= _GEN_285;
    end
    if (_T_440) begin
      _T_2304 <= 1'h0;
    end else begin
      _T_2304 <= _GEN_276;
    end
    if (_T_440) begin
      _T_2243 <= 1'h0;
    end else begin
      _T_2243 <= _GEN_267;
    end
    if (_T_440) begin
      _T_2182 <= 1'h0;
    end else begin
      _T_2182 <= _GEN_258;
    end
    if (_T_440) begin
      _T_2121 <= 1'h0;
    end else begin
      _T_2121 <= _GEN_249;
    end
    if (_T_440) begin
      _T_2060 <= 1'h0;
    end else begin
      _T_2060 <= _GEN_240;
    end
    if (_T_440) begin
      _T_1999 <= 1'h0;
    end else begin
      _T_1999 <= _GEN_231;
    end
    if (_T_440) begin
      _T_1938 <= 1'h0;
    end else begin
      _T_1938 <= _GEN_222;
    end
    if (_T_440) begin
      _T_1877 <= 1'h0;
    end else begin
      _T_1877 <= _GEN_213;
    end
    if (_T_440) begin
      _T_1816 <= 1'h0;
    end else begin
      _T_1816 <= _GEN_204;
    end
    if (_T_440) begin
      _T_1755 <= 1'h0;
    end else begin
      _T_1755 <= _GEN_195;
    end
    if (_T_440) begin
      _T_1694 <= 1'h0;
    end else begin
      _T_1694 <= _GEN_186;
    end
    if (_T_440) begin
      _T_1633 <= 1'h0;
    end else begin
      _T_1633 <= _GEN_177;
    end
    if (_T_440) begin
      _T_1572 <= 1'h0;
    end else begin
      _T_1572 <= _GEN_168;
    end
    if (_T_440) begin
      _T_1511 <= 1'h0;
    end else begin
      _T_1511 <= _GEN_159;
    end
    if (_T_440) begin
      _T_1450 <= 1'h0;
    end else begin
      _T_1450 <= _GEN_150;
    end
    if (_T_440) begin
      _T_1389 <= 1'h0;
    end else begin
      _T_1389 <= _GEN_141;
    end
    if (_T_440) begin
      _T_1328 <= 1'h0;
    end else begin
      _T_1328 <= _GEN_132;
    end
    if (_T_440) begin
      _T_1267 <= 1'h0;
    end else begin
      _T_1267 <= _GEN_123;
    end
    if (_T_440) begin
      _T_1206 <= 1'h0;
    end else begin
      _T_1206 <= _GEN_114;
    end
    if (_T_440) begin
      _T_1145 <= 1'h0;
    end else begin
      _T_1145 <= _GEN_105;
    end
    if (_T_440) begin
      _T_1084 <= 1'h0;
    end else begin
      _T_1084 <= _GEN_96;
    end
    if (_T_440) begin
      _T_1023 <= 1'h0;
    end else begin
      _T_1023 <= _GEN_87;
    end
    if (_T_440) begin
      _T_962 <= 1'h0;
    end else begin
      _T_962 <= _GEN_78;
    end
    if (_T_440) begin
      _T_901 <= 1'h0;
    end else begin
      _T_901 <= _GEN_69;
    end
    if (_T_440) begin
      _T_840 <= 1'h0;
    end else begin
      _T_840 <= _GEN_60;
    end
    if (_T_440) begin
      _T_779 <= 1'h0;
    end else begin
      _T_779 <= _GEN_51;
    end
    if (_T_440) begin
      _T_718 <= 1'h0;
    end else begin
      _T_718 <= _GEN_42;
    end
    if (_T_440) begin
      _T_657 <= 1'h0;
    end else begin
      _T_657 <= _GEN_33;
    end
    if (_T_440) begin
      _T_596 <= 1'h0;
    end else begin
      _T_596 <= _GEN_24;
    end
    if (_T_440) begin
      _T_535 <= 1'h0;
    end else begin
      _T_535 <= _GEN_15;
    end
    if (_T_440) begin
      _T_474 <= 1'h0;
    end else begin
      _T_474 <= _GEN_6;
    end
    if (reset) begin
      _T_4309 <= 22'h0;
    end else if (_T_4308) begin
      _T_4309 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4248 <= 22'h0;
    end else if (_T_4247) begin
      _T_4248 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4187 <= 22'h0;
    end else if (_T_4186) begin
      _T_4187 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4126 <= 22'h0;
    end else if (_T_4125) begin
      _T_4126 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4065 <= 22'h0;
    end else if (_T_4064) begin
      _T_4065 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4004 <= 22'h0;
    end else if (_T_4003) begin
      _T_4004 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3943 <= 22'h0;
    end else if (_T_3942) begin
      _T_3943 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3882 <= 22'h0;
    end else if (_T_3881) begin
      _T_3882 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3821 <= 22'h0;
    end else if (_T_3820) begin
      _T_3821 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3760 <= 22'h0;
    end else if (_T_3759) begin
      _T_3760 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3699 <= 22'h0;
    end else if (_T_3698) begin
      _T_3699 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3638 <= 22'h0;
    end else if (_T_3637) begin
      _T_3638 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3577 <= 22'h0;
    end else if (_T_3576) begin
      _T_3577 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3516 <= 22'h0;
    end else if (_T_3515) begin
      _T_3516 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3455 <= 22'h0;
    end else if (_T_3454) begin
      _T_3455 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3394 <= 22'h0;
    end else if (_T_3393) begin
      _T_3394 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3333 <= 22'h0;
    end else if (_T_3332) begin
      _T_3333 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3272 <= 22'h0;
    end else if (_T_3271) begin
      _T_3272 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3211 <= 22'h0;
    end else if (_T_3210) begin
      _T_3211 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3150 <= 22'h0;
    end else if (_T_3149) begin
      _T_3150 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3089 <= 22'h0;
    end else if (_T_3088) begin
      _T_3089 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3028 <= 22'h0;
    end else if (_T_3027) begin
      _T_3028 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2967 <= 22'h0;
    end else if (_T_2966) begin
      _T_2967 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2906 <= 22'h0;
    end else if (_T_2905) begin
      _T_2906 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2845 <= 22'h0;
    end else if (_T_2844) begin
      _T_2845 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2784 <= 22'h0;
    end else if (_T_2783) begin
      _T_2784 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2723 <= 22'h0;
    end else if (_T_2722) begin
      _T_2723 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2662 <= 22'h0;
    end else if (_T_2661) begin
      _T_2662 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2601 <= 22'h0;
    end else if (_T_2600) begin
      _T_2601 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2540 <= 22'h0;
    end else if (_T_2539) begin
      _T_2540 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2479 <= 22'h0;
    end else if (_T_2478) begin
      _T_2479 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2418 <= 22'h0;
    end else if (_T_2417) begin
      _T_2418 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2357 <= 22'h0;
    end else if (_T_2356) begin
      _T_2357 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2296 <= 22'h0;
    end else if (_T_2295) begin
      _T_2296 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2235 <= 22'h0;
    end else if (_T_2234) begin
      _T_2235 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2174 <= 22'h0;
    end else if (_T_2173) begin
      _T_2174 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2113 <= 22'h0;
    end else if (_T_2112) begin
      _T_2113 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2052 <= 22'h0;
    end else if (_T_2051) begin
      _T_2052 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1991 <= 22'h0;
    end else if (_T_1990) begin
      _T_1991 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1930 <= 22'h0;
    end else if (_T_1929) begin
      _T_1930 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1869 <= 22'h0;
    end else if (_T_1868) begin
      _T_1869 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1808 <= 22'h0;
    end else if (_T_1807) begin
      _T_1808 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1747 <= 22'h0;
    end else if (_T_1746) begin
      _T_1747 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1686 <= 22'h0;
    end else if (_T_1685) begin
      _T_1686 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1625 <= 22'h0;
    end else if (_T_1624) begin
      _T_1625 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1564 <= 22'h0;
    end else if (_T_1563) begin
      _T_1564 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1503 <= 22'h0;
    end else if (_T_1502) begin
      _T_1503 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1442 <= 22'h0;
    end else if (_T_1441) begin
      _T_1442 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1381 <= 22'h0;
    end else if (_T_1380) begin
      _T_1381 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1320 <= 22'h0;
    end else if (_T_1319) begin
      _T_1320 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1259 <= 22'h0;
    end else if (_T_1258) begin
      _T_1259 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1198 <= 22'h0;
    end else if (_T_1197) begin
      _T_1198 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1137 <= 22'h0;
    end else if (_T_1136) begin
      _T_1137 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1076 <= 22'h0;
    end else if (_T_1075) begin
      _T_1076 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1015 <= 22'h0;
    end else if (_T_1014) begin
      _T_1015 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_954 <= 22'h0;
    end else if (_T_953) begin
      _T_954 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_893 <= 22'h0;
    end else if (_T_892) begin
      _T_893 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_832 <= 22'h0;
    end else if (_T_831) begin
      _T_832 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_771 <= 22'h0;
    end else if (_T_770) begin
      _T_771 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_710 <= 22'h0;
    end else if (_T_709) begin
      _T_710 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_649 <= 22'h0;
    end else if (_T_648) begin
      _T_649 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_588 <= 22'h0;
    end else if (_T_587) begin
      _T_588 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_527 <= 22'h0;
    end else if (_T_526) begin
      _T_527 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_466 <= 22'h0;
    end else if (_T_465) begin
      _T_466 <= io_cacheIn_addr[31:10];
    end
    if (_T_440) begin
      _T_4331 <= 1'h0;
    end else begin
      _T_4331 <= _GEN_575;
    end
    if (_T_440) begin
      _T_4270 <= 1'h0;
    end else begin
      _T_4270 <= _GEN_566;
    end
    if (_T_440) begin
      _T_4209 <= 1'h0;
    end else begin
      _T_4209 <= _GEN_557;
    end
    if (_T_440) begin
      _T_4148 <= 1'h0;
    end else begin
      _T_4148 <= _GEN_548;
    end
    if (_T_440) begin
      _T_4087 <= 1'h0;
    end else begin
      _T_4087 <= _GEN_539;
    end
    if (_T_440) begin
      _T_4026 <= 1'h0;
    end else begin
      _T_4026 <= _GEN_530;
    end
    if (_T_440) begin
      _T_3965 <= 1'h0;
    end else begin
      _T_3965 <= _GEN_521;
    end
    if (_T_440) begin
      _T_3904 <= 1'h0;
    end else begin
      _T_3904 <= _GEN_512;
    end
    if (_T_440) begin
      _T_3843 <= 1'h0;
    end else begin
      _T_3843 <= _GEN_503;
    end
    if (_T_440) begin
      _T_3782 <= 1'h0;
    end else begin
      _T_3782 <= _GEN_494;
    end
    if (_T_440) begin
      _T_3721 <= 1'h0;
    end else begin
      _T_3721 <= _GEN_485;
    end
    if (_T_440) begin
      _T_3660 <= 1'h0;
    end else begin
      _T_3660 <= _GEN_476;
    end
    if (_T_440) begin
      _T_3599 <= 1'h0;
    end else begin
      _T_3599 <= _GEN_467;
    end
    if (_T_440) begin
      _T_3538 <= 1'h0;
    end else begin
      _T_3538 <= _GEN_458;
    end
    if (_T_440) begin
      _T_3477 <= 1'h0;
    end else begin
      _T_3477 <= _GEN_449;
    end
    if (_T_440) begin
      _T_3416 <= 1'h0;
    end else begin
      _T_3416 <= _GEN_440;
    end
    if (_T_440) begin
      _T_3355 <= 1'h0;
    end else begin
      _T_3355 <= _GEN_431;
    end
    if (_T_440) begin
      _T_3294 <= 1'h0;
    end else begin
      _T_3294 <= _GEN_422;
    end
    if (_T_440) begin
      _T_3233 <= 1'h0;
    end else begin
      _T_3233 <= _GEN_413;
    end
    if (_T_440) begin
      _T_3172 <= 1'h0;
    end else begin
      _T_3172 <= _GEN_404;
    end
    if (_T_440) begin
      _T_3111 <= 1'h0;
    end else begin
      _T_3111 <= _GEN_395;
    end
    if (_T_440) begin
      _T_3050 <= 1'h0;
    end else begin
      _T_3050 <= _GEN_386;
    end
    if (_T_440) begin
      _T_2989 <= 1'h0;
    end else begin
      _T_2989 <= _GEN_377;
    end
    if (_T_440) begin
      _T_2928 <= 1'h0;
    end else begin
      _T_2928 <= _GEN_368;
    end
    if (_T_440) begin
      _T_2867 <= 1'h0;
    end else begin
      _T_2867 <= _GEN_359;
    end
    if (_T_440) begin
      _T_2806 <= 1'h0;
    end else begin
      _T_2806 <= _GEN_350;
    end
    if (_T_440) begin
      _T_2745 <= 1'h0;
    end else begin
      _T_2745 <= _GEN_341;
    end
    if (_T_440) begin
      _T_2684 <= 1'h0;
    end else begin
      _T_2684 <= _GEN_332;
    end
    if (_T_440) begin
      _T_2623 <= 1'h0;
    end else begin
      _T_2623 <= _GEN_323;
    end
    if (_T_440) begin
      _T_2562 <= 1'h0;
    end else begin
      _T_2562 <= _GEN_314;
    end
    if (_T_440) begin
      _T_2501 <= 1'h0;
    end else begin
      _T_2501 <= _GEN_305;
    end
    if (_T_440) begin
      _T_2440 <= 1'h0;
    end else begin
      _T_2440 <= _GEN_296;
    end
    if (_T_440) begin
      _T_2379 <= 1'h0;
    end else begin
      _T_2379 <= _GEN_287;
    end
    if (_T_440) begin
      _T_2318 <= 1'h0;
    end else begin
      _T_2318 <= _GEN_278;
    end
    if (_T_440) begin
      _T_2257 <= 1'h0;
    end else begin
      _T_2257 <= _GEN_269;
    end
    if (_T_440) begin
      _T_2196 <= 1'h0;
    end else begin
      _T_2196 <= _GEN_260;
    end
    if (_T_440) begin
      _T_2135 <= 1'h0;
    end else begin
      _T_2135 <= _GEN_251;
    end
    if (_T_440) begin
      _T_2074 <= 1'h0;
    end else begin
      _T_2074 <= _GEN_242;
    end
    if (_T_440) begin
      _T_2013 <= 1'h0;
    end else begin
      _T_2013 <= _GEN_233;
    end
    if (_T_440) begin
      _T_1952 <= 1'h0;
    end else begin
      _T_1952 <= _GEN_224;
    end
    if (_T_440) begin
      _T_1891 <= 1'h0;
    end else begin
      _T_1891 <= _GEN_215;
    end
    if (_T_440) begin
      _T_1830 <= 1'h0;
    end else begin
      _T_1830 <= _GEN_206;
    end
    if (_T_440) begin
      _T_1769 <= 1'h0;
    end else begin
      _T_1769 <= _GEN_197;
    end
    if (_T_440) begin
      _T_1708 <= 1'h0;
    end else begin
      _T_1708 <= _GEN_188;
    end
    if (_T_440) begin
      _T_1647 <= 1'h0;
    end else begin
      _T_1647 <= _GEN_179;
    end
    if (_T_440) begin
      _T_1586 <= 1'h0;
    end else begin
      _T_1586 <= _GEN_170;
    end
    if (_T_440) begin
      _T_1525 <= 1'h0;
    end else begin
      _T_1525 <= _GEN_161;
    end
    if (_T_440) begin
      _T_1464 <= 1'h0;
    end else begin
      _T_1464 <= _GEN_152;
    end
    if (_T_440) begin
      _T_1403 <= 1'h0;
    end else begin
      _T_1403 <= _GEN_143;
    end
    if (_T_440) begin
      _T_1342 <= 1'h0;
    end else begin
      _T_1342 <= _GEN_134;
    end
    if (_T_440) begin
      _T_1281 <= 1'h0;
    end else begin
      _T_1281 <= _GEN_125;
    end
    if (_T_440) begin
      _T_1220 <= 1'h0;
    end else begin
      _T_1220 <= _GEN_116;
    end
    if (_T_440) begin
      _T_1159 <= 1'h0;
    end else begin
      _T_1159 <= _GEN_107;
    end
    if (_T_440) begin
      _T_1098 <= 1'h0;
    end else begin
      _T_1098 <= _GEN_98;
    end
    if (_T_440) begin
      _T_1037 <= 1'h0;
    end else begin
      _T_1037 <= _GEN_89;
    end
    if (_T_440) begin
      _T_976 <= 1'h0;
    end else begin
      _T_976 <= _GEN_80;
    end
    if (_T_440) begin
      _T_915 <= 1'h0;
    end else begin
      _T_915 <= _GEN_71;
    end
    if (_T_440) begin
      _T_854 <= 1'h0;
    end else begin
      _T_854 <= _GEN_62;
    end
    if (_T_440) begin
      _T_793 <= 1'h0;
    end else begin
      _T_793 <= _GEN_53;
    end
    if (_T_440) begin
      _T_732 <= 1'h0;
    end else begin
      _T_732 <= _GEN_44;
    end
    if (_T_440) begin
      _T_671 <= 1'h0;
    end else begin
      _T_671 <= _GEN_35;
    end
    if (_T_440) begin
      _T_610 <= 1'h0;
    end else begin
      _T_610 <= _GEN_26;
    end
    if (_T_440) begin
      _T_549 <= 1'h0;
    end else begin
      _T_549 <= _GEN_17;
    end
    if (_T_440) begin
      _T_488 <= 1'h0;
    end else begin
      _T_488 <= _GEN_8;
    end
    if (reset) begin
      _T_4323 <= 22'h0;
    end else if (_T_4322) begin
      _T_4323 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4262 <= 22'h0;
    end else if (_T_4261) begin
      _T_4262 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4201 <= 22'h0;
    end else if (_T_4200) begin
      _T_4201 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4140 <= 22'h0;
    end else if (_T_4139) begin
      _T_4140 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4079 <= 22'h0;
    end else if (_T_4078) begin
      _T_4079 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4018 <= 22'h0;
    end else if (_T_4017) begin
      _T_4018 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3957 <= 22'h0;
    end else if (_T_3956) begin
      _T_3957 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3896 <= 22'h0;
    end else if (_T_3895) begin
      _T_3896 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3835 <= 22'h0;
    end else if (_T_3834) begin
      _T_3835 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3774 <= 22'h0;
    end else if (_T_3773) begin
      _T_3774 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3713 <= 22'h0;
    end else if (_T_3712) begin
      _T_3713 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3652 <= 22'h0;
    end else if (_T_3651) begin
      _T_3652 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3591 <= 22'h0;
    end else if (_T_3590) begin
      _T_3591 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3530 <= 22'h0;
    end else if (_T_3529) begin
      _T_3530 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3469 <= 22'h0;
    end else if (_T_3468) begin
      _T_3469 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3408 <= 22'h0;
    end else if (_T_3407) begin
      _T_3408 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3347 <= 22'h0;
    end else if (_T_3346) begin
      _T_3347 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3286 <= 22'h0;
    end else if (_T_3285) begin
      _T_3286 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3225 <= 22'h0;
    end else if (_T_3224) begin
      _T_3225 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3164 <= 22'h0;
    end else if (_T_3163) begin
      _T_3164 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3103 <= 22'h0;
    end else if (_T_3102) begin
      _T_3103 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3042 <= 22'h0;
    end else if (_T_3041) begin
      _T_3042 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2981 <= 22'h0;
    end else if (_T_2980) begin
      _T_2981 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2920 <= 22'h0;
    end else if (_T_2919) begin
      _T_2920 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2859 <= 22'h0;
    end else if (_T_2858) begin
      _T_2859 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2798 <= 22'h0;
    end else if (_T_2797) begin
      _T_2798 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2737 <= 22'h0;
    end else if (_T_2736) begin
      _T_2737 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2676 <= 22'h0;
    end else if (_T_2675) begin
      _T_2676 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2615 <= 22'h0;
    end else if (_T_2614) begin
      _T_2615 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2554 <= 22'h0;
    end else if (_T_2553) begin
      _T_2554 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2493 <= 22'h0;
    end else if (_T_2492) begin
      _T_2493 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2432 <= 22'h0;
    end else if (_T_2431) begin
      _T_2432 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2371 <= 22'h0;
    end else if (_T_2370) begin
      _T_2371 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2310 <= 22'h0;
    end else if (_T_2309) begin
      _T_2310 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2249 <= 22'h0;
    end else if (_T_2248) begin
      _T_2249 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2188 <= 22'h0;
    end else if (_T_2187) begin
      _T_2188 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2127 <= 22'h0;
    end else if (_T_2126) begin
      _T_2127 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2066 <= 22'h0;
    end else if (_T_2065) begin
      _T_2066 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2005 <= 22'h0;
    end else if (_T_2004) begin
      _T_2005 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1944 <= 22'h0;
    end else if (_T_1943) begin
      _T_1944 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1883 <= 22'h0;
    end else if (_T_1882) begin
      _T_1883 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1822 <= 22'h0;
    end else if (_T_1821) begin
      _T_1822 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1761 <= 22'h0;
    end else if (_T_1760) begin
      _T_1761 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1700 <= 22'h0;
    end else if (_T_1699) begin
      _T_1700 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1639 <= 22'h0;
    end else if (_T_1638) begin
      _T_1639 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1578 <= 22'h0;
    end else if (_T_1577) begin
      _T_1578 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1517 <= 22'h0;
    end else if (_T_1516) begin
      _T_1517 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1456 <= 22'h0;
    end else if (_T_1455) begin
      _T_1456 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1395 <= 22'h0;
    end else if (_T_1394) begin
      _T_1395 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1334 <= 22'h0;
    end else if (_T_1333) begin
      _T_1334 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1273 <= 22'h0;
    end else if (_T_1272) begin
      _T_1273 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1212 <= 22'h0;
    end else if (_T_1211) begin
      _T_1212 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1151 <= 22'h0;
    end else if (_T_1150) begin
      _T_1151 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1090 <= 22'h0;
    end else if (_T_1089) begin
      _T_1090 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1029 <= 22'h0;
    end else if (_T_1028) begin
      _T_1029 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_968 <= 22'h0;
    end else if (_T_967) begin
      _T_968 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_907 <= 22'h0;
    end else if (_T_906) begin
      _T_907 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_846 <= 22'h0;
    end else if (_T_845) begin
      _T_846 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_785 <= 22'h0;
    end else if (_T_784) begin
      _T_785 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_724 <= 22'h0;
    end else if (_T_723) begin
      _T_724 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_663 <= 22'h0;
    end else if (_T_662) begin
      _T_663 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_602 <= 22'h0;
    end else if (_T_601) begin
      _T_602 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_541 <= 22'h0;
    end else if (_T_540) begin
      _T_541 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_480 <= 22'h0;
    end else if (_T_479) begin
      _T_480 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_493 <= 2'h0;
    end else if (_T_492) begin
      _T_493 <= _T_490;
    end
    if (reset) begin
      _T_432 <= 2'h0;
    end else if (_T_431) begin
      _T_432 <= _T_429;
    end
    if (reset) begin
      _T_554 <= 2'h0;
    end else if (_T_553) begin
      _T_554 <= _T_551;
    end
    if (reset) begin
      _T_615 <= 2'h0;
    end else if (_T_614) begin
      _T_615 <= _T_612;
    end
    if (reset) begin
      _T_676 <= 2'h0;
    end else if (_T_675) begin
      _T_676 <= _T_673;
    end
    if (reset) begin
      _T_737 <= 2'h0;
    end else if (_T_736) begin
      _T_737 <= _T_734;
    end
    if (reset) begin
      _T_798 <= 2'h0;
    end else if (_T_797) begin
      _T_798 <= _T_795;
    end
    if (reset) begin
      _T_859 <= 2'h0;
    end else if (_T_858) begin
      _T_859 <= _T_856;
    end
    if (reset) begin
      _T_920 <= 2'h0;
    end else if (_T_919) begin
      _T_920 <= _T_917;
    end
    if (reset) begin
      _T_981 <= 2'h0;
    end else if (_T_980) begin
      _T_981 <= _T_978;
    end
    if (reset) begin
      _T_1042 <= 2'h0;
    end else if (_T_1041) begin
      _T_1042 <= _T_1039;
    end
    if (reset) begin
      _T_1103 <= 2'h0;
    end else if (_T_1102) begin
      _T_1103 <= _T_1100;
    end
    if (reset) begin
      _T_1164 <= 2'h0;
    end else if (_T_1163) begin
      _T_1164 <= _T_1161;
    end
    if (reset) begin
      _T_1225 <= 2'h0;
    end else if (_T_1224) begin
      _T_1225 <= _T_1222;
    end
    if (reset) begin
      _T_1286 <= 2'h0;
    end else if (_T_1285) begin
      _T_1286 <= _T_1283;
    end
    if (reset) begin
      _T_1347 <= 2'h0;
    end else if (_T_1346) begin
      _T_1347 <= _T_1344;
    end
    if (reset) begin
      _T_1408 <= 2'h0;
    end else if (_T_1407) begin
      _T_1408 <= _T_1405;
    end
    if (reset) begin
      _T_1469 <= 2'h0;
    end else if (_T_1468) begin
      _T_1469 <= _T_1466;
    end
    if (reset) begin
      _T_1530 <= 2'h0;
    end else if (_T_1529) begin
      _T_1530 <= _T_1527;
    end
    if (reset) begin
      _T_1591 <= 2'h0;
    end else if (_T_1590) begin
      _T_1591 <= _T_1588;
    end
    if (reset) begin
      _T_1652 <= 2'h0;
    end else if (_T_1651) begin
      _T_1652 <= _T_1649;
    end
    if (reset) begin
      _T_1713 <= 2'h0;
    end else if (_T_1712) begin
      _T_1713 <= _T_1710;
    end
    if (reset) begin
      _T_1774 <= 2'h0;
    end else if (_T_1773) begin
      _T_1774 <= _T_1771;
    end
    if (reset) begin
      _T_1835 <= 2'h0;
    end else if (_T_1834) begin
      _T_1835 <= _T_1832;
    end
    if (reset) begin
      _T_1896 <= 2'h0;
    end else if (_T_1895) begin
      _T_1896 <= _T_1893;
    end
    if (reset) begin
      _T_1957 <= 2'h0;
    end else if (_T_1956) begin
      _T_1957 <= _T_1954;
    end
    if (reset) begin
      _T_2018 <= 2'h0;
    end else if (_T_2017) begin
      _T_2018 <= _T_2015;
    end
    if (reset) begin
      _T_2079 <= 2'h0;
    end else if (_T_2078) begin
      _T_2079 <= _T_2076;
    end
    if (reset) begin
      _T_2140 <= 2'h0;
    end else if (_T_2139) begin
      _T_2140 <= _T_2137;
    end
    if (reset) begin
      _T_2201 <= 2'h0;
    end else if (_T_2200) begin
      _T_2201 <= _T_2198;
    end
    if (reset) begin
      _T_2262 <= 2'h0;
    end else if (_T_2261) begin
      _T_2262 <= _T_2259;
    end
    if (reset) begin
      _T_2323 <= 2'h0;
    end else if (_T_2322) begin
      _T_2323 <= _T_2320;
    end
    if (reset) begin
      _T_2384 <= 2'h0;
    end else if (_T_2383) begin
      _T_2384 <= _T_2381;
    end
    if (reset) begin
      _T_2445 <= 2'h0;
    end else if (_T_2444) begin
      _T_2445 <= _T_2442;
    end
    if (reset) begin
      _T_2506 <= 2'h0;
    end else if (_T_2505) begin
      _T_2506 <= _T_2503;
    end
    if (reset) begin
      _T_2567 <= 2'h0;
    end else if (_T_2566) begin
      _T_2567 <= _T_2564;
    end
    if (reset) begin
      _T_2628 <= 2'h0;
    end else if (_T_2627) begin
      _T_2628 <= _T_2625;
    end
    if (reset) begin
      _T_2689 <= 2'h0;
    end else if (_T_2688) begin
      _T_2689 <= _T_2686;
    end
    if (reset) begin
      _T_2750 <= 2'h0;
    end else if (_T_2749) begin
      _T_2750 <= _T_2747;
    end
    if (reset) begin
      _T_2811 <= 2'h0;
    end else if (_T_2810) begin
      _T_2811 <= _T_2808;
    end
    if (reset) begin
      _T_2872 <= 2'h0;
    end else if (_T_2871) begin
      _T_2872 <= _T_2869;
    end
    if (reset) begin
      _T_2933 <= 2'h0;
    end else if (_T_2932) begin
      _T_2933 <= _T_2930;
    end
    if (reset) begin
      _T_2994 <= 2'h0;
    end else if (_T_2993) begin
      _T_2994 <= _T_2991;
    end
    if (reset) begin
      _T_3055 <= 2'h0;
    end else if (_T_3054) begin
      _T_3055 <= _T_3052;
    end
    if (reset) begin
      _T_3116 <= 2'h0;
    end else if (_T_3115) begin
      _T_3116 <= _T_3113;
    end
    if (reset) begin
      _T_3177 <= 2'h0;
    end else if (_T_3176) begin
      _T_3177 <= _T_3174;
    end
    if (reset) begin
      _T_3238 <= 2'h0;
    end else if (_T_3237) begin
      _T_3238 <= _T_3235;
    end
    if (reset) begin
      _T_3299 <= 2'h0;
    end else if (_T_3298) begin
      _T_3299 <= _T_3296;
    end
    if (reset) begin
      _T_3360 <= 2'h0;
    end else if (_T_3359) begin
      _T_3360 <= _T_3357;
    end
    if (reset) begin
      _T_3421 <= 2'h0;
    end else if (_T_3420) begin
      _T_3421 <= _T_3418;
    end
    if (reset) begin
      _T_3482 <= 2'h0;
    end else if (_T_3481) begin
      _T_3482 <= _T_3479;
    end
    if (reset) begin
      _T_3543 <= 2'h0;
    end else if (_T_3542) begin
      _T_3543 <= _T_3540;
    end
    if (reset) begin
      _T_3604 <= 2'h0;
    end else if (_T_3603) begin
      _T_3604 <= _T_3601;
    end
    if (reset) begin
      _T_3665 <= 2'h0;
    end else if (_T_3664) begin
      _T_3665 <= _T_3662;
    end
    if (reset) begin
      _T_3726 <= 2'h0;
    end else if (_T_3725) begin
      _T_3726 <= _T_3723;
    end
    if (reset) begin
      _T_3787 <= 2'h0;
    end else if (_T_3786) begin
      _T_3787 <= _T_3784;
    end
    if (reset) begin
      _T_3848 <= 2'h0;
    end else if (_T_3847) begin
      _T_3848 <= _T_3845;
    end
    if (reset) begin
      _T_3909 <= 2'h0;
    end else if (_T_3908) begin
      _T_3909 <= _T_3906;
    end
    if (reset) begin
      _T_3970 <= 2'h0;
    end else if (_T_3969) begin
      _T_3970 <= _T_3967;
    end
    if (reset) begin
      _T_4031 <= 2'h0;
    end else if (_T_4030) begin
      _T_4031 <= _T_4028;
    end
    if (reset) begin
      _T_4092 <= 2'h0;
    end else if (_T_4091) begin
      _T_4092 <= _T_4089;
    end
    if (reset) begin
      _T_4153 <= 2'h0;
    end else if (_T_4152) begin
      _T_4153 <= _T_4150;
    end
    if (reset) begin
      _T_4214 <= 2'h0;
    end else if (_T_4213) begin
      _T_4214 <= _T_4211;
    end
    if (reset) begin
      _T_4275 <= 2'h0;
    end else if (_T_4274) begin
      _T_4275 <= _T_4272;
    end
  end
endmodule
module AXICache(
  input         clock,
  input         reset,
  input         io_axiIO_awready,
  output        io_axiIO_awvalid,
  output [31:0] io_axiIO_awaddr,
  output [2:0]  io_axiIO_awsize,
  input         io_axiIO_wready,
  output        io_axiIO_wvalid,
  output [63:0] io_axiIO_wdata,
  output [7:0]  io_axiIO_wstrb,
  output        io_axiIO_wlast,
  output        io_axiIO_bready,
  input         io_axiIO_bvalid,
  input         io_axiIO_arready,
  output        io_axiIO_arvalid,
  output [31:0] io_axiIO_araddr,
  output [7:0]  io_axiIO_arlen,
  output [2:0]  io_axiIO_arsize,
  output [1:0]  io_axiIO_arburst,
  output        io_axiIO_rready,
  input         io_axiIO_rvalid,
  input  [63:0] io_axiIO_rdata,
  input         io_axiIO_rlast,
  input         io_cache_ar_valid_o,
  input  [31:0] io_cache_ar_addr_o,
  input  [7:0]  io_cache_ar_len_o,
  output        io_cache_r_valid_i,
  output [63:0] io_cache_r_data_i,
  output        io_cache_r_last_i,
  input         io_cache_w_valid_o,
  output        io_cache_w_ready_i,
  input  [63:0] io_cache_w_data_o,
  input  [31:0] io_cache_w_addr_o,
  input  [7:0]  io_cache_w_mask_o,
  input  [1:0]  io_cache_wsize
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] rd_state; // @[AXICache.scala 26:25]
  wire  _T = io_axiIO_rlast & io_axiIO_rvalid; // @[AXICache.scala 31:22]
  wire  _T_3 = 2'h0 == rd_state; // @[Mux.scala 80:60]
  wire  _T_5 = 2'h1 == rd_state; // @[Mux.scala 80:60]
  wire  _T_7 = 2'h2 == rd_state; // @[Mux.scala 80:60]
  wire  isReq = rd_state == 2'h1; // @[AXICache.scala 47:24]
  wire  isData = rd_state == 2'h2; // @[AXICache.scala 48:25]
  wire [1:0] _T_12 = isReq ? 2'h3 : 2'h0; // @[AXICache.scala 63:25]
  wire [1:0] valid_c = {io_axiIO_awready,io_axiIO_wready}; // @[Cat.scala 29:58]
  reg [1:0] w_state; // @[AXICache.scala 76:24]
  wire  _T_15 = 2'h2 == valid_c; // @[Mux.scala 80:60]
  wire  _T_17 = 2'h3 == valid_c; // @[Mux.scala 80:60]
  wire  _T_18 = 2'h1 == w_state; // @[Mux.scala 80:60]
  wire  _T_20 = 2'h2 == w_state; // @[Mux.scala 80:60]
  wire  _T_22 = 2'h3 == w_state; // @[Mux.scala 80:60]
  wire  isWReq = w_state == 2'h1; // @[AXICache.scala 100:24]
  wire  isWData = w_state == 2'h2; // @[AXICache.scala 101:25]
  wire  isWB = w_state == 2'h3; // @[AXICache.scala 102:22]
  wire  _T_27 = isWReq | isWData; // @[AXICache.scala 127:29]
  assign io_axiIO_awvalid = w_state == 2'h1; // @[AXICache.scala 118:20]
  assign io_axiIO_awaddr = isWReq ? io_cache_w_addr_o : 32'h0; // @[AXICache.scala 119:19]
  assign io_axiIO_awsize = {{1'd0}, io_cache_wsize}; // @[AXICache.scala 122:19]
  assign io_axiIO_wvalid = isWReq | isWData; // @[AXICache.scala 127:19]
  assign io_axiIO_wdata = _T_27 ? io_cache_w_data_o : 64'h0; // @[AXICache.scala 128:18]
  assign io_axiIO_wstrb = _T_27 ? io_cache_w_mask_o : 8'h0; // @[AXICache.scala 129:18]
  assign io_axiIO_wlast = isWReq | isWData; // @[AXICache.scala 130:18]
  assign io_axiIO_bready = w_state == 2'h3; // @[AXICache.scala 133:19]
  assign io_axiIO_arvalid = rd_state == 2'h1; // @[AXICache.scala 59:19]
  assign io_axiIO_araddr = isReq ? io_cache_ar_addr_o : 32'h0; // @[AXICache.scala 60:19]
  assign io_axiIO_arlen = isReq ? io_cache_ar_len_o : 8'h0; // @[AXICache.scala 62:18]
  assign io_axiIO_arsize = {{1'd0}, _T_12}; // @[AXICache.scala 63:19]
  assign io_axiIO_arburst = isReq ? 2'h1 : 2'h0; // @[AXICache.scala 64:20]
  assign io_axiIO_rready = isData | isReq; // @[AXICache.scala 67:18]
  assign io_cache_r_valid_i = io_axiIO_rvalid; // @[AXICache.scala 52:22]
  assign io_cache_r_data_i = io_axiIO_rdata; // @[AXICache.scala 53:21]
  assign io_cache_r_last_i = io_axiIO_rlast; // @[AXICache.scala 51:21]
  assign io_cache_w_ready_i = io_axiIO_bvalid & isWB; // @[AXICache.scala 104:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rd_state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  w_state = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      rd_state <= 2'h0;
    end else if (_T_7) begin
      if (_T) begin
        rd_state <= 2'h0;
      end else begin
        rd_state <= 2'h2;
      end
    end else if (_T_5) begin
      if (io_axiIO_arready) begin
        if (_T) begin
          rd_state <= 2'h0;
        end else begin
          rd_state <= 2'h2;
        end
      end else begin
        rd_state <= 2'h1;
      end
    end else if (_T_3) begin
      if (io_cache_ar_valid_o) begin
        rd_state <= 2'h1;
      end else begin
        rd_state <= 2'h0;
      end
    end
    if (reset) begin
      w_state <= 2'h0;
    end else if (_T_22) begin
      if (io_axiIO_bvalid) begin
        w_state <= 2'h0;
      end else begin
        w_state <= 2'h3;
      end
    end else if (_T_20) begin
      if (io_axiIO_wready) begin
        w_state <= 2'h3;
      end else begin
        w_state <= 2'h2;
      end
    end else if (_T_18) begin
      if (_T_17) begin
        w_state <= 2'h3;
      end else if (_T_15) begin
        w_state <= 2'h2;
      end else begin
        w_state <= 2'h1;
      end
    end else if (io_cache_w_valid_o) begin
      w_state <= 2'h1;
    end else begin
      w_state <= 2'h0;
    end
  end
endmodule
module arbTop(
  input         io_arbIn_valid,
  output        io_arbIn_ready,
  output [63:0] io_arbIn_data_read,
  input  [63:0] io_arbIn_data_write,
  input         io_arbIn_wen,
  input  [31:0] io_arbIn_addr,
  input  [1:0]  io_arbIn_rsize,
  input  [7:0]  io_arbIn_mask,
  output        io_arbMMIO_valid,
  input         io_arbMMIO_ready,
  input  [63:0] io_arbMMIO_data_read,
  output [63:0] io_arbMMIO_data_write,
  output        io_arbMMIO_wen,
  output [31:0] io_arbMMIO_addr,
  output [1:0]  io_arbMMIO_rsize,
  output [7:0]  io_arbMMIO_mask,
  output        io_arbClint_valid,
  input  [63:0] io_arbClint_data_read,
  output [63:0] io_arbClint_data_write,
  output        io_arbClint_wen,
  output [31:0] io_arbClint_addr,
  output        io_arbDCache_valid,
  input         io_arbDCache_ready,
  input  [63:0] io_arbDCache_data_read,
  output [63:0] io_arbDCache_data_write,
  output        io_arbDCache_wen,
  output [31:0] io_arbDCache_addr,
  output [1:0]  io_arbDCache_rsize,
  output [7:0]  io_arbDCache_mask,
  output        io_arbCgra_valid,
  input         io_arbCgra_ready,
  input  [63:0] io_arbCgra_data_read,
  output [63:0] io_arbCgra_data_write,
  output        io_arbCgra_wen,
  output [31:0] io_arbCgra_addr
);
  wire  _T = io_arbIn_addr >= 32'h2000000; // @[arbCpu2Cache.scala 153:31]
  wire  _T_1 = io_arbIn_addr < 32'h200bfff; // @[arbCpu2Cache.scala 153:61]
  wire  clinitV = _T & _T_1; // @[arbCpu2Cache.scala 153:45]
  wire  _T_2 = io_arbIn_addr >= 32'h80000000; // @[arbCpu2Cache.scala 154:31]
  wire  _T_3 = io_arbIn_addr < 32'h8fffffff; // @[arbCpu2Cache.scala 154:60]
  wire  dCacheV = _T_2 & _T_3; // @[arbCpu2Cache.scala 154:44]
  wire  mmioV = io_arbIn_addr >= 32'h8fffffff; // @[arbCpu2Cache.scala 155:29]
  wire  _T_7 = ~clinitV; // @[arbCpu2Cache.scala 160:25]
  wire  _T_8 = ~dCacheV; // @[arbCpu2Cache.scala 160:37]
  wire  _T_9 = _T_7 & _T_8; // @[arbCpu2Cache.scala 160:34]
  wire  _T_10 = ~mmioV; // @[arbCpu2Cache.scala 160:49]
  wire  _T_11 = _T_9 & _T_10; // @[arbCpu2Cache.scala 160:46]
  wire  _T_14 = dCacheV & io_arbDCache_ready; // @[arbCpu2Cache.scala 170:63]
  wire  _T_15 = clinitV | _T_14; // @[arbCpu2Cache.scala 170:51]
  wire  _T_16 = mmioV & io_arbMMIO_ready; // @[arbCpu2Cache.scala 170:96]
  wire  _T_17 = _T_15 | _T_16; // @[arbCpu2Cache.scala 170:86]
  wire  _T_23 = _T_11 & io_arbCgra_ready; // @[arbCpu2Cache.scala 170:153]
  wire [63:0] _T_25 = mmioV ? io_arbMMIO_data_read : io_arbCgra_data_read; // @[arbCpu2Cache.scala 171:97]
  wire [63:0] _T_26 = clinitV ? io_arbClint_data_read : _T_25; // @[arbCpu2Cache.scala 171:63]
  assign io_arbIn_ready = _T_17 | _T_23; // @[arbCpu2Cache.scala 170:18]
  assign io_arbIn_data_read = dCacheV ? io_arbDCache_data_read : _T_26; // @[arbCpu2Cache.scala 171:22]
  assign io_arbMMIO_valid = mmioV & io_arbIn_valid; // @[arbCpu2Cache.scala 159:20]
  assign io_arbMMIO_data_write = io_arbIn_data_write; // @[arbCpu2Cache.scala 163:23]
  assign io_arbMMIO_wen = io_arbIn_wen; // @[arbCpu2Cache.scala 163:23]
  assign io_arbMMIO_addr = io_arbIn_addr; // @[arbCpu2Cache.scala 163:23]
  assign io_arbMMIO_rsize = io_arbIn_rsize; // @[arbCpu2Cache.scala 163:23]
  assign io_arbMMIO_mask = io_arbIn_mask; // @[arbCpu2Cache.scala 163:23]
  assign io_arbClint_valid = clinitV & io_arbIn_valid; // @[arbCpu2Cache.scala 157:21]
  assign io_arbClint_data_write = io_arbIn_data_write; // @[arbCpu2Cache.scala 164:24]
  assign io_arbClint_wen = io_arbIn_wen; // @[arbCpu2Cache.scala 164:24]
  assign io_arbClint_addr = io_arbIn_addr; // @[arbCpu2Cache.scala 164:24]
  assign io_arbDCache_valid = dCacheV & io_arbIn_valid; // @[arbCpu2Cache.scala 158:22]
  assign io_arbDCache_data_write = io_arbIn_data_write; // @[arbCpu2Cache.scala 165:25]
  assign io_arbDCache_wen = io_arbIn_wen; // @[arbCpu2Cache.scala 165:25]
  assign io_arbDCache_addr = io_arbIn_addr; // @[arbCpu2Cache.scala 165:25]
  assign io_arbDCache_rsize = io_arbIn_rsize; // @[arbCpu2Cache.scala 165:25]
  assign io_arbDCache_mask = io_arbIn_mask; // @[arbCpu2Cache.scala 165:25]
  assign io_arbCgra_valid = _T_11 & io_arbIn_valid; // @[arbCpu2Cache.scala 160:20]
  assign io_arbCgra_data_write = io_arbIn_data_write; // @[arbCpu2Cache.scala 166:23]
  assign io_arbCgra_wen = io_arbIn_wen; // @[arbCpu2Cache.scala 166:23]
  assign io_arbCgra_addr = io_arbIn_addr; // @[arbCpu2Cache.scala 166:23]
endmodule
module mmioCache(
  input         io_mmioIn_valid,
  output        io_mmioIn_ready,
  output [63:0] io_mmioIn_data_read,
  input  [63:0] io_mmioIn_data_write,
  input         io_mmioIn_wen,
  input  [31:0] io_mmioIn_addr,
  output        io_mmioOut_valid,
  input         io_mmioOut_ready,
  input  [63:0] io_mmioOut_data_read,
  output [63:0] io_mmioOut_data_write,
  output        io_mmioOut_wen,
  output [31:0] io_mmioOut_addr
);
  assign io_mmioIn_ready = io_mmioOut_ready; // @[mmioCache.scala 14:12]
  assign io_mmioIn_data_read = io_mmioOut_data_read; // @[mmioCache.scala 14:12]
  assign io_mmioOut_valid = io_mmioIn_valid; // @[mmioCache.scala 14:12]
  assign io_mmioOut_data_write = io_mmioIn_data_write; // @[mmioCache.scala 14:12]
  assign io_mmioOut_wen = io_mmioIn_wen; // @[mmioCache.scala 14:12]
  assign io_mmioOut_addr = io_mmioIn_addr; // @[mmioCache.scala 14:12]
endmodule
module Dcache(
  input          clock,
  input          reset,
  output         io_cacheOut_ar_valid_o,
  output [31:0]  io_cacheOut_ar_addr_o,
  output [7:0]   io_cacheOut_ar_len_o,
  input          io_cacheOut_r_valid_i,
  input  [63:0]  io_cacheOut_r_data_i,
  input          io_cacheOut_r_last_i,
  output         io_cacheOut_w_valid_o,
  input          io_cacheOut_w_ready_i,
  output [63:0]  io_cacheOut_w_data_o,
  output [31:0]  io_cacheOut_w_addr_o,
  output [7:0]   io_cacheOut_w_mask_o,
  output [1:0]   io_cacheOut_wsize,
  input          io_cacheIn_valid,
  output         io_cacheIn_ready,
  output [63:0]  io_cacheIn_data_read,
  input  [63:0]  io_cacheIn_data_write,
  input          io_cacheIn_wen,
  input  [31:0]  io_cacheIn_addr,
  input  [1:0]   io_cacheIn_rsize,
  input  [7:0]   io_cacheIn_mask,
  output         io_SRAMIO_0_cen,
  output         io_SRAMIO_0_wen,
  output [127:0] io_SRAMIO_0_wdata,
  output [5:0]   io_SRAMIO_0_addr,
  output [127:0] io_SRAMIO_0_wmask,
  input  [127:0] io_SRAMIO_0_rdata,
  output         io_SRAMIO_1_cen,
  output         io_SRAMIO_1_wen,
  output [127:0] io_SRAMIO_1_wdata,
  output [5:0]   io_SRAMIO_1_addr,
  output [127:0] io_SRAMIO_1_wmask,
  input  [127:0] io_SRAMIO_1_rdata,
  output         io_SRAMIO_2_cen,
  output         io_SRAMIO_2_wen,
  output [127:0] io_SRAMIO_2_wdata,
  output [5:0]   io_SRAMIO_2_addr,
  output [127:0] io_SRAMIO_2_wmask,
  input  [127:0] io_SRAMIO_2_rdata,
  output         io_SRAMIO_3_cen,
  output         io_SRAMIO_3_wen,
  output [127:0] io_SRAMIO_3_wdata,
  output [5:0]   io_SRAMIO_3_addr,
  output [127:0] io_SRAMIO_3_wmask,
  input  [127:0] io_SRAMIO_3_rdata,
  input          io_block,
  input          updataICache
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] _T_4; // @[Cache.scala 704:29]
  wire  _T_281 = 6'h3f == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_4297; // @[Reg.scala 27:20]
  wire  _T_279 = 6'h3e == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_4236; // @[Reg.scala 27:20]
  wire  _T_277 = 6'h3d == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_4175; // @[Reg.scala 27:20]
  wire  _T_275 = 6'h3c == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_4114; // @[Reg.scala 27:20]
  wire  _T_273 = 6'h3b == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_4053; // @[Reg.scala 27:20]
  wire  _T_271 = 6'h3a == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3992; // @[Reg.scala 27:20]
  wire  _T_269 = 6'h39 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3931; // @[Reg.scala 27:20]
  wire  _T_267 = 6'h38 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3870; // @[Reg.scala 27:20]
  wire  _T_265 = 6'h37 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3809; // @[Reg.scala 27:20]
  wire  _T_263 = 6'h36 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3748; // @[Reg.scala 27:20]
  wire  _T_261 = 6'h35 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3687; // @[Reg.scala 27:20]
  wire  _T_259 = 6'h34 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3626; // @[Reg.scala 27:20]
  wire  _T_257 = 6'h33 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3565; // @[Reg.scala 27:20]
  wire  _T_255 = 6'h32 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3504; // @[Reg.scala 27:20]
  wire  _T_253 = 6'h31 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3443; // @[Reg.scala 27:20]
  wire  _T_251 = 6'h30 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3382; // @[Reg.scala 27:20]
  wire  _T_249 = 6'h2f == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3321; // @[Reg.scala 27:20]
  wire  _T_247 = 6'h2e == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3260; // @[Reg.scala 27:20]
  wire  _T_245 = 6'h2d == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3199; // @[Reg.scala 27:20]
  wire  _T_243 = 6'h2c == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3138; // @[Reg.scala 27:20]
  wire  _T_241 = 6'h2b == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3077; // @[Reg.scala 27:20]
  wire  _T_239 = 6'h2a == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_3016; // @[Reg.scala 27:20]
  wire  _T_237 = 6'h29 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2955; // @[Reg.scala 27:20]
  wire  _T_235 = 6'h28 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2894; // @[Reg.scala 27:20]
  wire  _T_233 = 6'h27 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2833; // @[Reg.scala 27:20]
  wire  _T_231 = 6'h26 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2772; // @[Reg.scala 27:20]
  wire  _T_229 = 6'h25 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2711; // @[Reg.scala 27:20]
  wire  _T_227 = 6'h24 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2650; // @[Reg.scala 27:20]
  wire  _T_225 = 6'h23 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2589; // @[Reg.scala 27:20]
  wire  _T_223 = 6'h22 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2528; // @[Reg.scala 27:20]
  wire  _T_221 = 6'h21 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2467; // @[Reg.scala 27:20]
  wire  _T_219 = 6'h20 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2406; // @[Reg.scala 27:20]
  wire  _T_217 = 6'h1f == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2345; // @[Reg.scala 27:20]
  wire  _T_215 = 6'h1e == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2284; // @[Reg.scala 27:20]
  wire  _T_213 = 6'h1d == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2223; // @[Reg.scala 27:20]
  wire  _T_211 = 6'h1c == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2162; // @[Reg.scala 27:20]
  wire  _T_209 = 6'h1b == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2101; // @[Reg.scala 27:20]
  wire  _T_207 = 6'h1a == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_2040; // @[Reg.scala 27:20]
  wire  _T_205 = 6'h19 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1979; // @[Reg.scala 27:20]
  wire  _T_203 = 6'h18 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1918; // @[Reg.scala 27:20]
  wire  _T_201 = 6'h17 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1857; // @[Reg.scala 27:20]
  wire  _T_199 = 6'h16 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1796; // @[Reg.scala 27:20]
  wire  _T_197 = 6'h15 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1735; // @[Reg.scala 27:20]
  wire  _T_195 = 6'h14 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1674; // @[Reg.scala 27:20]
  wire  _T_193 = 6'h13 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1613; // @[Reg.scala 27:20]
  wire  _T_191 = 6'h12 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1552; // @[Reg.scala 27:20]
  wire  _T_189 = 6'h11 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1491; // @[Reg.scala 27:20]
  wire  _T_187 = 6'h10 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1430; // @[Reg.scala 27:20]
  wire  _T_185 = 6'hf == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1369; // @[Reg.scala 27:20]
  wire  _T_183 = 6'he == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1308; // @[Reg.scala 27:20]
  wire  _T_181 = 6'hd == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1247; // @[Reg.scala 27:20]
  wire  _T_179 = 6'hc == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1186; // @[Reg.scala 27:20]
  wire  _T_177 = 6'hb == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1125; // @[Reg.scala 27:20]
  wire  _T_175 = 6'ha == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1064; // @[Reg.scala 27:20]
  wire  _T_173 = 6'h9 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_1003; // @[Reg.scala 27:20]
  wire  _T_171 = 6'h8 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_942; // @[Reg.scala 27:20]
  wire  _T_169 = 6'h7 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_881; // @[Reg.scala 27:20]
  wire  _T_167 = 6'h6 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_820; // @[Reg.scala 27:20]
  wire  _T_165 = 6'h5 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_759; // @[Reg.scala 27:20]
  wire  _T_163 = 6'h4 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_698; // @[Reg.scala 27:20]
  wire  _T_161 = 6'h3 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_637; // @[Reg.scala 27:20]
  wire  _T_159 = 6'h2 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_576; // @[Reg.scala 27:20]
  wire  _T_157 = 6'h1 == io_cacheIn_addr[9:4]; // @[Mux.scala 80:60]
  reg  _T_515; // @[Reg.scala 27:20]
  reg  _T_454; // @[Reg.scala 27:20]
  wire  _T_158_0 = _T_157 ? _T_515 : _T_454; // @[Mux.scala 80:57]
  wire  _T_160_0 = _T_159 ? _T_576 : _T_158_0; // @[Mux.scala 80:57]
  wire  _T_162_0 = _T_161 ? _T_637 : _T_160_0; // @[Mux.scala 80:57]
  wire  _T_164_0 = _T_163 ? _T_698 : _T_162_0; // @[Mux.scala 80:57]
  wire  _T_166_0 = _T_165 ? _T_759 : _T_164_0; // @[Mux.scala 80:57]
  wire  _T_168_0 = _T_167 ? _T_820 : _T_166_0; // @[Mux.scala 80:57]
  wire  _T_170_0 = _T_169 ? _T_881 : _T_168_0; // @[Mux.scala 80:57]
  wire  _T_172_0 = _T_171 ? _T_942 : _T_170_0; // @[Mux.scala 80:57]
  wire  _T_174_0 = _T_173 ? _T_1003 : _T_172_0; // @[Mux.scala 80:57]
  wire  _T_176_0 = _T_175 ? _T_1064 : _T_174_0; // @[Mux.scala 80:57]
  wire  _T_178_0 = _T_177 ? _T_1125 : _T_176_0; // @[Mux.scala 80:57]
  wire  _T_180_0 = _T_179 ? _T_1186 : _T_178_0; // @[Mux.scala 80:57]
  wire  _T_182_0 = _T_181 ? _T_1247 : _T_180_0; // @[Mux.scala 80:57]
  wire  _T_184_0 = _T_183 ? _T_1308 : _T_182_0; // @[Mux.scala 80:57]
  wire  _T_186_0 = _T_185 ? _T_1369 : _T_184_0; // @[Mux.scala 80:57]
  wire  _T_188_0 = _T_187 ? _T_1430 : _T_186_0; // @[Mux.scala 80:57]
  wire  _T_190_0 = _T_189 ? _T_1491 : _T_188_0; // @[Mux.scala 80:57]
  wire  _T_192_0 = _T_191 ? _T_1552 : _T_190_0; // @[Mux.scala 80:57]
  wire  _T_194_0 = _T_193 ? _T_1613 : _T_192_0; // @[Mux.scala 80:57]
  wire  _T_196_0 = _T_195 ? _T_1674 : _T_194_0; // @[Mux.scala 80:57]
  wire  _T_198_0 = _T_197 ? _T_1735 : _T_196_0; // @[Mux.scala 80:57]
  wire  _T_200_0 = _T_199 ? _T_1796 : _T_198_0; // @[Mux.scala 80:57]
  wire  _T_202_0 = _T_201 ? _T_1857 : _T_200_0; // @[Mux.scala 80:57]
  wire  _T_204_0 = _T_203 ? _T_1918 : _T_202_0; // @[Mux.scala 80:57]
  wire  _T_206_0 = _T_205 ? _T_1979 : _T_204_0; // @[Mux.scala 80:57]
  wire  _T_208_0 = _T_207 ? _T_2040 : _T_206_0; // @[Mux.scala 80:57]
  wire  _T_210_0 = _T_209 ? _T_2101 : _T_208_0; // @[Mux.scala 80:57]
  wire  _T_212_0 = _T_211 ? _T_2162 : _T_210_0; // @[Mux.scala 80:57]
  wire  _T_214_0 = _T_213 ? _T_2223 : _T_212_0; // @[Mux.scala 80:57]
  wire  _T_216_0 = _T_215 ? _T_2284 : _T_214_0; // @[Mux.scala 80:57]
  wire  _T_218_0 = _T_217 ? _T_2345 : _T_216_0; // @[Mux.scala 80:57]
  wire  _T_220_0 = _T_219 ? _T_2406 : _T_218_0; // @[Mux.scala 80:57]
  wire  _T_222_0 = _T_221 ? _T_2467 : _T_220_0; // @[Mux.scala 80:57]
  wire  _T_224_0 = _T_223 ? _T_2528 : _T_222_0; // @[Mux.scala 80:57]
  wire  _T_226_0 = _T_225 ? _T_2589 : _T_224_0; // @[Mux.scala 80:57]
  wire  _T_228_0 = _T_227 ? _T_2650 : _T_226_0; // @[Mux.scala 80:57]
  wire  _T_230_0 = _T_229 ? _T_2711 : _T_228_0; // @[Mux.scala 80:57]
  wire  _T_232_0 = _T_231 ? _T_2772 : _T_230_0; // @[Mux.scala 80:57]
  wire  _T_234_0 = _T_233 ? _T_2833 : _T_232_0; // @[Mux.scala 80:57]
  wire  _T_236_0 = _T_235 ? _T_2894 : _T_234_0; // @[Mux.scala 80:57]
  wire  _T_238_0 = _T_237 ? _T_2955 : _T_236_0; // @[Mux.scala 80:57]
  wire  _T_240_0 = _T_239 ? _T_3016 : _T_238_0; // @[Mux.scala 80:57]
  wire  _T_242_0 = _T_241 ? _T_3077 : _T_240_0; // @[Mux.scala 80:57]
  wire  _T_244_0 = _T_243 ? _T_3138 : _T_242_0; // @[Mux.scala 80:57]
  wire  _T_246_0 = _T_245 ? _T_3199 : _T_244_0; // @[Mux.scala 80:57]
  wire  _T_248_0 = _T_247 ? _T_3260 : _T_246_0; // @[Mux.scala 80:57]
  wire  _T_250_0 = _T_249 ? _T_3321 : _T_248_0; // @[Mux.scala 80:57]
  wire  _T_252_0 = _T_251 ? _T_3382 : _T_250_0; // @[Mux.scala 80:57]
  wire  _T_254_0 = _T_253 ? _T_3443 : _T_252_0; // @[Mux.scala 80:57]
  wire  _T_256_0 = _T_255 ? _T_3504 : _T_254_0; // @[Mux.scala 80:57]
  wire  _T_258_0 = _T_257 ? _T_3565 : _T_256_0; // @[Mux.scala 80:57]
  wire  _T_260_0 = _T_259 ? _T_3626 : _T_258_0; // @[Mux.scala 80:57]
  wire  _T_262_0 = _T_261 ? _T_3687 : _T_260_0; // @[Mux.scala 80:57]
  wire  _T_264_0 = _T_263 ? _T_3748 : _T_262_0; // @[Mux.scala 80:57]
  wire  _T_266_0 = _T_265 ? _T_3809 : _T_264_0; // @[Mux.scala 80:57]
  wire  _T_268_0 = _T_267 ? _T_3870 : _T_266_0; // @[Mux.scala 80:57]
  wire  _T_270_0 = _T_269 ? _T_3931 : _T_268_0; // @[Mux.scala 80:57]
  wire  _T_272_0 = _T_271 ? _T_3992 : _T_270_0; // @[Mux.scala 80:57]
  wire  _T_274_0 = _T_273 ? _T_4053 : _T_272_0; // @[Mux.scala 80:57]
  wire  _T_276_0 = _T_275 ? _T_4114 : _T_274_0; // @[Mux.scala 80:57]
  wire  _T_278_0 = _T_277 ? _T_4175 : _T_276_0; // @[Mux.scala 80:57]
  wire  _T_280_0 = _T_279 ? _T_4236 : _T_278_0; // @[Mux.scala 80:57]
  wire  _T_282_0 = _T_281 ? _T_4297 : _T_280_0; // @[Mux.scala 80:57]
  reg [21:0] _T_4289; // @[Reg.scala 27:20]
  reg [21:0] _T_4228; // @[Reg.scala 27:20]
  reg [21:0] _T_4167; // @[Reg.scala 27:20]
  reg [21:0] _T_4106; // @[Reg.scala 27:20]
  reg [21:0] _T_4045; // @[Reg.scala 27:20]
  reg [21:0] _T_3984; // @[Reg.scala 27:20]
  reg [21:0] _T_3923; // @[Reg.scala 27:20]
  reg [21:0] _T_3862; // @[Reg.scala 27:20]
  reg [21:0] _T_3801; // @[Reg.scala 27:20]
  reg [21:0] _T_3740; // @[Reg.scala 27:20]
  reg [21:0] _T_3679; // @[Reg.scala 27:20]
  reg [21:0] _T_3618; // @[Reg.scala 27:20]
  reg [21:0] _T_3557; // @[Reg.scala 27:20]
  reg [21:0] _T_3496; // @[Reg.scala 27:20]
  reg [21:0] _T_3435; // @[Reg.scala 27:20]
  reg [21:0] _T_3374; // @[Reg.scala 27:20]
  reg [21:0] _T_3313; // @[Reg.scala 27:20]
  reg [21:0] _T_3252; // @[Reg.scala 27:20]
  reg [21:0] _T_3191; // @[Reg.scala 27:20]
  reg [21:0] _T_3130; // @[Reg.scala 27:20]
  reg [21:0] _T_3069; // @[Reg.scala 27:20]
  reg [21:0] _T_3008; // @[Reg.scala 27:20]
  reg [21:0] _T_2947; // @[Reg.scala 27:20]
  reg [21:0] _T_2886; // @[Reg.scala 27:20]
  reg [21:0] _T_2825; // @[Reg.scala 27:20]
  reg [21:0] _T_2764; // @[Reg.scala 27:20]
  reg [21:0] _T_2703; // @[Reg.scala 27:20]
  reg [21:0] _T_2642; // @[Reg.scala 27:20]
  reg [21:0] _T_2581; // @[Reg.scala 27:20]
  reg [21:0] _T_2520; // @[Reg.scala 27:20]
  reg [21:0] _T_2459; // @[Reg.scala 27:20]
  reg [21:0] _T_2398; // @[Reg.scala 27:20]
  reg [21:0] _T_2337; // @[Reg.scala 27:20]
  reg [21:0] _T_2276; // @[Reg.scala 27:20]
  reg [21:0] _T_2215; // @[Reg.scala 27:20]
  reg [21:0] _T_2154; // @[Reg.scala 27:20]
  reg [21:0] _T_2093; // @[Reg.scala 27:20]
  reg [21:0] _T_2032; // @[Reg.scala 27:20]
  reg [21:0] _T_1971; // @[Reg.scala 27:20]
  reg [21:0] _T_1910; // @[Reg.scala 27:20]
  reg [21:0] _T_1849; // @[Reg.scala 27:20]
  reg [21:0] _T_1788; // @[Reg.scala 27:20]
  reg [21:0] _T_1727; // @[Reg.scala 27:20]
  reg [21:0] _T_1666; // @[Reg.scala 27:20]
  reg [21:0] _T_1605; // @[Reg.scala 27:20]
  reg [21:0] _T_1544; // @[Reg.scala 27:20]
  reg [21:0] _T_1483; // @[Reg.scala 27:20]
  reg [21:0] _T_1422; // @[Reg.scala 27:20]
  reg [21:0] _T_1361; // @[Reg.scala 27:20]
  reg [21:0] _T_1300; // @[Reg.scala 27:20]
  reg [21:0] _T_1239; // @[Reg.scala 27:20]
  reg [21:0] _T_1178; // @[Reg.scala 27:20]
  reg [21:0] _T_1117; // @[Reg.scala 27:20]
  reg [21:0] _T_1056; // @[Reg.scala 27:20]
  reg [21:0] _T_995; // @[Reg.scala 27:20]
  reg [21:0] _T_934; // @[Reg.scala 27:20]
  reg [21:0] _T_873; // @[Reg.scala 27:20]
  reg [21:0] _T_812; // @[Reg.scala 27:20]
  reg [21:0] _T_751; // @[Reg.scala 27:20]
  reg [21:0] _T_690; // @[Reg.scala 27:20]
  reg [21:0] _T_629; // @[Reg.scala 27:20]
  reg [21:0] _T_568; // @[Reg.scala 27:20]
  reg [21:0] _T_507; // @[Reg.scala 27:20]
  reg [21:0] _T_446; // @[Reg.scala 27:20]
  wire [21:0] _T_32_0 = _T_157 ? _T_507 : _T_446; // @[Mux.scala 80:57]
  wire [21:0] _T_34_0 = _T_159 ? _T_568 : _T_32_0; // @[Mux.scala 80:57]
  wire [21:0] _T_36_0 = _T_161 ? _T_629 : _T_34_0; // @[Mux.scala 80:57]
  wire [21:0] _T_38_0 = _T_163 ? _T_690 : _T_36_0; // @[Mux.scala 80:57]
  wire [21:0] _T_40_0 = _T_165 ? _T_751 : _T_38_0; // @[Mux.scala 80:57]
  wire [21:0] _T_42_0 = _T_167 ? _T_812 : _T_40_0; // @[Mux.scala 80:57]
  wire [21:0] _T_44_0 = _T_169 ? _T_873 : _T_42_0; // @[Mux.scala 80:57]
  wire [21:0] _T_46_0 = _T_171 ? _T_934 : _T_44_0; // @[Mux.scala 80:57]
  wire [21:0] _T_48_0 = _T_173 ? _T_995 : _T_46_0; // @[Mux.scala 80:57]
  wire [21:0] _T_50_0 = _T_175 ? _T_1056 : _T_48_0; // @[Mux.scala 80:57]
  wire [21:0] _T_52_0 = _T_177 ? _T_1117 : _T_50_0; // @[Mux.scala 80:57]
  wire [21:0] _T_54_0 = _T_179 ? _T_1178 : _T_52_0; // @[Mux.scala 80:57]
  wire [21:0] _T_56_0 = _T_181 ? _T_1239 : _T_54_0; // @[Mux.scala 80:57]
  wire [21:0] _T_58_0 = _T_183 ? _T_1300 : _T_56_0; // @[Mux.scala 80:57]
  wire [21:0] _T_60_0 = _T_185 ? _T_1361 : _T_58_0; // @[Mux.scala 80:57]
  wire [21:0] _T_62_0 = _T_187 ? _T_1422 : _T_60_0; // @[Mux.scala 80:57]
  wire [21:0] _T_64_0 = _T_189 ? _T_1483 : _T_62_0; // @[Mux.scala 80:57]
  wire [21:0] _T_66_0 = _T_191 ? _T_1544 : _T_64_0; // @[Mux.scala 80:57]
  wire [21:0] _T_68_0 = _T_193 ? _T_1605 : _T_66_0; // @[Mux.scala 80:57]
  wire [21:0] _T_70_0 = _T_195 ? _T_1666 : _T_68_0; // @[Mux.scala 80:57]
  wire [21:0] _T_72_0 = _T_197 ? _T_1727 : _T_70_0; // @[Mux.scala 80:57]
  wire [21:0] _T_74_0 = _T_199 ? _T_1788 : _T_72_0; // @[Mux.scala 80:57]
  wire [21:0] _T_76_0 = _T_201 ? _T_1849 : _T_74_0; // @[Mux.scala 80:57]
  wire [21:0] _T_78_0 = _T_203 ? _T_1910 : _T_76_0; // @[Mux.scala 80:57]
  wire [21:0] _T_80_0 = _T_205 ? _T_1971 : _T_78_0; // @[Mux.scala 80:57]
  wire [21:0] _T_82_0 = _T_207 ? _T_2032 : _T_80_0; // @[Mux.scala 80:57]
  wire [21:0] _T_84_0 = _T_209 ? _T_2093 : _T_82_0; // @[Mux.scala 80:57]
  wire [21:0] _T_86_0 = _T_211 ? _T_2154 : _T_84_0; // @[Mux.scala 80:57]
  wire [21:0] _T_88_0 = _T_213 ? _T_2215 : _T_86_0; // @[Mux.scala 80:57]
  wire [21:0] _T_90_0 = _T_215 ? _T_2276 : _T_88_0; // @[Mux.scala 80:57]
  wire [21:0] _T_92_0 = _T_217 ? _T_2337 : _T_90_0; // @[Mux.scala 80:57]
  wire [21:0] _T_94_0 = _T_219 ? _T_2398 : _T_92_0; // @[Mux.scala 80:57]
  wire [21:0] _T_96_0 = _T_221 ? _T_2459 : _T_94_0; // @[Mux.scala 80:57]
  wire [21:0] _T_98_0 = _T_223 ? _T_2520 : _T_96_0; // @[Mux.scala 80:57]
  wire [21:0] _T_100_0 = _T_225 ? _T_2581 : _T_98_0; // @[Mux.scala 80:57]
  wire [21:0] _T_102_0 = _T_227 ? _T_2642 : _T_100_0; // @[Mux.scala 80:57]
  wire [21:0] _T_104_0 = _T_229 ? _T_2703 : _T_102_0; // @[Mux.scala 80:57]
  wire [21:0] _T_106_0 = _T_231 ? _T_2764 : _T_104_0; // @[Mux.scala 80:57]
  wire [21:0] _T_108_0 = _T_233 ? _T_2825 : _T_106_0; // @[Mux.scala 80:57]
  wire [21:0] _T_110_0 = _T_235 ? _T_2886 : _T_108_0; // @[Mux.scala 80:57]
  wire [21:0] _T_112_0 = _T_237 ? _T_2947 : _T_110_0; // @[Mux.scala 80:57]
  wire [21:0] _T_114_0 = _T_239 ? _T_3008 : _T_112_0; // @[Mux.scala 80:57]
  wire [21:0] _T_116_0 = _T_241 ? _T_3069 : _T_114_0; // @[Mux.scala 80:57]
  wire [21:0] _T_118_0 = _T_243 ? _T_3130 : _T_116_0; // @[Mux.scala 80:57]
  wire [21:0] _T_120_0 = _T_245 ? _T_3191 : _T_118_0; // @[Mux.scala 80:57]
  wire [21:0] _T_122_0 = _T_247 ? _T_3252 : _T_120_0; // @[Mux.scala 80:57]
  wire [21:0] _T_124_0 = _T_249 ? _T_3313 : _T_122_0; // @[Mux.scala 80:57]
  wire [21:0] _T_126_0 = _T_251 ? _T_3374 : _T_124_0; // @[Mux.scala 80:57]
  wire [21:0] _T_128_0 = _T_253 ? _T_3435 : _T_126_0; // @[Mux.scala 80:57]
  wire [21:0] _T_130_0 = _T_255 ? _T_3496 : _T_128_0; // @[Mux.scala 80:57]
  wire [21:0] _T_132_0 = _T_257 ? _T_3557 : _T_130_0; // @[Mux.scala 80:57]
  wire [21:0] _T_134_0 = _T_259 ? _T_3618 : _T_132_0; // @[Mux.scala 80:57]
  wire [21:0] _T_136_0 = _T_261 ? _T_3679 : _T_134_0; // @[Mux.scala 80:57]
  wire [21:0] _T_138_0 = _T_263 ? _T_3740 : _T_136_0; // @[Mux.scala 80:57]
  wire [21:0] _T_140_0 = _T_265 ? _T_3801 : _T_138_0; // @[Mux.scala 80:57]
  wire [21:0] _T_142_0 = _T_267 ? _T_3862 : _T_140_0; // @[Mux.scala 80:57]
  wire [21:0] _T_144_0 = _T_269 ? _T_3923 : _T_142_0; // @[Mux.scala 80:57]
  wire [21:0] _T_146_0 = _T_271 ? _T_3984 : _T_144_0; // @[Mux.scala 80:57]
  wire [21:0] _T_148_0 = _T_273 ? _T_4045 : _T_146_0; // @[Mux.scala 80:57]
  wire [21:0] _T_150_0 = _T_275 ? _T_4106 : _T_148_0; // @[Mux.scala 80:57]
  wire [21:0] _T_152_0 = _T_277 ? _T_4167 : _T_150_0; // @[Mux.scala 80:57]
  wire [21:0] _T_154_0 = _T_279 ? _T_4228 : _T_152_0; // @[Mux.scala 80:57]
  wire [21:0] _T_156_0 = _T_281 ? _T_4289 : _T_154_0; // @[Mux.scala 80:57]
  wire  _T_283 = _T_156_0 == io_cacheIn_addr[31:10]; // @[Cache.scala 772:78]
  wire  _T_284 = _T_282_0 & _T_283; // @[Cache.scala 772:62]
  reg  _T_4311; // @[Reg.scala 27:20]
  reg  _T_4250; // @[Reg.scala 27:20]
  reg  _T_4189; // @[Reg.scala 27:20]
  reg  _T_4128; // @[Reg.scala 27:20]
  reg  _T_4067; // @[Reg.scala 27:20]
  reg  _T_4006; // @[Reg.scala 27:20]
  reg  _T_3945; // @[Reg.scala 27:20]
  reg  _T_3884; // @[Reg.scala 27:20]
  reg  _T_3823; // @[Reg.scala 27:20]
  reg  _T_3762; // @[Reg.scala 27:20]
  reg  _T_3701; // @[Reg.scala 27:20]
  reg  _T_3640; // @[Reg.scala 27:20]
  reg  _T_3579; // @[Reg.scala 27:20]
  reg  _T_3518; // @[Reg.scala 27:20]
  reg  _T_3457; // @[Reg.scala 27:20]
  reg  _T_3396; // @[Reg.scala 27:20]
  reg  _T_3335; // @[Reg.scala 27:20]
  reg  _T_3274; // @[Reg.scala 27:20]
  reg  _T_3213; // @[Reg.scala 27:20]
  reg  _T_3152; // @[Reg.scala 27:20]
  reg  _T_3091; // @[Reg.scala 27:20]
  reg  _T_3030; // @[Reg.scala 27:20]
  reg  _T_2969; // @[Reg.scala 27:20]
  reg  _T_2908; // @[Reg.scala 27:20]
  reg  _T_2847; // @[Reg.scala 27:20]
  reg  _T_2786; // @[Reg.scala 27:20]
  reg  _T_2725; // @[Reg.scala 27:20]
  reg  _T_2664; // @[Reg.scala 27:20]
  reg  _T_2603; // @[Reg.scala 27:20]
  reg  _T_2542; // @[Reg.scala 27:20]
  reg  _T_2481; // @[Reg.scala 27:20]
  reg  _T_2420; // @[Reg.scala 27:20]
  reg  _T_2359; // @[Reg.scala 27:20]
  reg  _T_2298; // @[Reg.scala 27:20]
  reg  _T_2237; // @[Reg.scala 27:20]
  reg  _T_2176; // @[Reg.scala 27:20]
  reg  _T_2115; // @[Reg.scala 27:20]
  reg  _T_2054; // @[Reg.scala 27:20]
  reg  _T_1993; // @[Reg.scala 27:20]
  reg  _T_1932; // @[Reg.scala 27:20]
  reg  _T_1871; // @[Reg.scala 27:20]
  reg  _T_1810; // @[Reg.scala 27:20]
  reg  _T_1749; // @[Reg.scala 27:20]
  reg  _T_1688; // @[Reg.scala 27:20]
  reg  _T_1627; // @[Reg.scala 27:20]
  reg  _T_1566; // @[Reg.scala 27:20]
  reg  _T_1505; // @[Reg.scala 27:20]
  reg  _T_1444; // @[Reg.scala 27:20]
  reg  _T_1383; // @[Reg.scala 27:20]
  reg  _T_1322; // @[Reg.scala 27:20]
  reg  _T_1261; // @[Reg.scala 27:20]
  reg  _T_1200; // @[Reg.scala 27:20]
  reg  _T_1139; // @[Reg.scala 27:20]
  reg  _T_1078; // @[Reg.scala 27:20]
  reg  _T_1017; // @[Reg.scala 27:20]
  reg  _T_956; // @[Reg.scala 27:20]
  reg  _T_895; // @[Reg.scala 27:20]
  reg  _T_834; // @[Reg.scala 27:20]
  reg  _T_773; // @[Reg.scala 27:20]
  reg  _T_712; // @[Reg.scala 27:20]
  reg  _T_651; // @[Reg.scala 27:20]
  reg  _T_590; // @[Reg.scala 27:20]
  reg  _T_529; // @[Reg.scala 27:20]
  reg  _T_468; // @[Reg.scala 27:20]
  wire  _T_158_1 = _T_157 ? _T_529 : _T_468; // @[Mux.scala 80:57]
  wire  _T_160_1 = _T_159 ? _T_590 : _T_158_1; // @[Mux.scala 80:57]
  wire  _T_162_1 = _T_161 ? _T_651 : _T_160_1; // @[Mux.scala 80:57]
  wire  _T_164_1 = _T_163 ? _T_712 : _T_162_1; // @[Mux.scala 80:57]
  wire  _T_166_1 = _T_165 ? _T_773 : _T_164_1; // @[Mux.scala 80:57]
  wire  _T_168_1 = _T_167 ? _T_834 : _T_166_1; // @[Mux.scala 80:57]
  wire  _T_170_1 = _T_169 ? _T_895 : _T_168_1; // @[Mux.scala 80:57]
  wire  _T_172_1 = _T_171 ? _T_956 : _T_170_1; // @[Mux.scala 80:57]
  wire  _T_174_1 = _T_173 ? _T_1017 : _T_172_1; // @[Mux.scala 80:57]
  wire  _T_176_1 = _T_175 ? _T_1078 : _T_174_1; // @[Mux.scala 80:57]
  wire  _T_178_1 = _T_177 ? _T_1139 : _T_176_1; // @[Mux.scala 80:57]
  wire  _T_180_1 = _T_179 ? _T_1200 : _T_178_1; // @[Mux.scala 80:57]
  wire  _T_182_1 = _T_181 ? _T_1261 : _T_180_1; // @[Mux.scala 80:57]
  wire  _T_184_1 = _T_183 ? _T_1322 : _T_182_1; // @[Mux.scala 80:57]
  wire  _T_186_1 = _T_185 ? _T_1383 : _T_184_1; // @[Mux.scala 80:57]
  wire  _T_188_1 = _T_187 ? _T_1444 : _T_186_1; // @[Mux.scala 80:57]
  wire  _T_190_1 = _T_189 ? _T_1505 : _T_188_1; // @[Mux.scala 80:57]
  wire  _T_192_1 = _T_191 ? _T_1566 : _T_190_1; // @[Mux.scala 80:57]
  wire  _T_194_1 = _T_193 ? _T_1627 : _T_192_1; // @[Mux.scala 80:57]
  wire  _T_196_1 = _T_195 ? _T_1688 : _T_194_1; // @[Mux.scala 80:57]
  wire  _T_198_1 = _T_197 ? _T_1749 : _T_196_1; // @[Mux.scala 80:57]
  wire  _T_200_1 = _T_199 ? _T_1810 : _T_198_1; // @[Mux.scala 80:57]
  wire  _T_202_1 = _T_201 ? _T_1871 : _T_200_1; // @[Mux.scala 80:57]
  wire  _T_204_1 = _T_203 ? _T_1932 : _T_202_1; // @[Mux.scala 80:57]
  wire  _T_206_1 = _T_205 ? _T_1993 : _T_204_1; // @[Mux.scala 80:57]
  wire  _T_208_1 = _T_207 ? _T_2054 : _T_206_1; // @[Mux.scala 80:57]
  wire  _T_210_1 = _T_209 ? _T_2115 : _T_208_1; // @[Mux.scala 80:57]
  wire  _T_212_1 = _T_211 ? _T_2176 : _T_210_1; // @[Mux.scala 80:57]
  wire  _T_214_1 = _T_213 ? _T_2237 : _T_212_1; // @[Mux.scala 80:57]
  wire  _T_216_1 = _T_215 ? _T_2298 : _T_214_1; // @[Mux.scala 80:57]
  wire  _T_218_1 = _T_217 ? _T_2359 : _T_216_1; // @[Mux.scala 80:57]
  wire  _T_220_1 = _T_219 ? _T_2420 : _T_218_1; // @[Mux.scala 80:57]
  wire  _T_222_1 = _T_221 ? _T_2481 : _T_220_1; // @[Mux.scala 80:57]
  wire  _T_224_1 = _T_223 ? _T_2542 : _T_222_1; // @[Mux.scala 80:57]
  wire  _T_226_1 = _T_225 ? _T_2603 : _T_224_1; // @[Mux.scala 80:57]
  wire  _T_228_1 = _T_227 ? _T_2664 : _T_226_1; // @[Mux.scala 80:57]
  wire  _T_230_1 = _T_229 ? _T_2725 : _T_228_1; // @[Mux.scala 80:57]
  wire  _T_232_1 = _T_231 ? _T_2786 : _T_230_1; // @[Mux.scala 80:57]
  wire  _T_234_1 = _T_233 ? _T_2847 : _T_232_1; // @[Mux.scala 80:57]
  wire  _T_236_1 = _T_235 ? _T_2908 : _T_234_1; // @[Mux.scala 80:57]
  wire  _T_238_1 = _T_237 ? _T_2969 : _T_236_1; // @[Mux.scala 80:57]
  wire  _T_240_1 = _T_239 ? _T_3030 : _T_238_1; // @[Mux.scala 80:57]
  wire  _T_242_1 = _T_241 ? _T_3091 : _T_240_1; // @[Mux.scala 80:57]
  wire  _T_244_1 = _T_243 ? _T_3152 : _T_242_1; // @[Mux.scala 80:57]
  wire  _T_246_1 = _T_245 ? _T_3213 : _T_244_1; // @[Mux.scala 80:57]
  wire  _T_248_1 = _T_247 ? _T_3274 : _T_246_1; // @[Mux.scala 80:57]
  wire  _T_250_1 = _T_249 ? _T_3335 : _T_248_1; // @[Mux.scala 80:57]
  wire  _T_252_1 = _T_251 ? _T_3396 : _T_250_1; // @[Mux.scala 80:57]
  wire  _T_254_1 = _T_253 ? _T_3457 : _T_252_1; // @[Mux.scala 80:57]
  wire  _T_256_1 = _T_255 ? _T_3518 : _T_254_1; // @[Mux.scala 80:57]
  wire  _T_258_1 = _T_257 ? _T_3579 : _T_256_1; // @[Mux.scala 80:57]
  wire  _T_260_1 = _T_259 ? _T_3640 : _T_258_1; // @[Mux.scala 80:57]
  wire  _T_262_1 = _T_261 ? _T_3701 : _T_260_1; // @[Mux.scala 80:57]
  wire  _T_264_1 = _T_263 ? _T_3762 : _T_262_1; // @[Mux.scala 80:57]
  wire  _T_266_1 = _T_265 ? _T_3823 : _T_264_1; // @[Mux.scala 80:57]
  wire  _T_268_1 = _T_267 ? _T_3884 : _T_266_1; // @[Mux.scala 80:57]
  wire  _T_270_1 = _T_269 ? _T_3945 : _T_268_1; // @[Mux.scala 80:57]
  wire  _T_272_1 = _T_271 ? _T_4006 : _T_270_1; // @[Mux.scala 80:57]
  wire  _T_274_1 = _T_273 ? _T_4067 : _T_272_1; // @[Mux.scala 80:57]
  wire  _T_276_1 = _T_275 ? _T_4128 : _T_274_1; // @[Mux.scala 80:57]
  wire  _T_278_1 = _T_277 ? _T_4189 : _T_276_1; // @[Mux.scala 80:57]
  wire  _T_280_1 = _T_279 ? _T_4250 : _T_278_1; // @[Mux.scala 80:57]
  wire  _T_282_1 = _T_281 ? _T_4311 : _T_280_1; // @[Mux.scala 80:57]
  reg [21:0] _T_4303; // @[Reg.scala 27:20]
  reg [21:0] _T_4242; // @[Reg.scala 27:20]
  reg [21:0] _T_4181; // @[Reg.scala 27:20]
  reg [21:0] _T_4120; // @[Reg.scala 27:20]
  reg [21:0] _T_4059; // @[Reg.scala 27:20]
  reg [21:0] _T_3998; // @[Reg.scala 27:20]
  reg [21:0] _T_3937; // @[Reg.scala 27:20]
  reg [21:0] _T_3876; // @[Reg.scala 27:20]
  reg [21:0] _T_3815; // @[Reg.scala 27:20]
  reg [21:0] _T_3754; // @[Reg.scala 27:20]
  reg [21:0] _T_3693; // @[Reg.scala 27:20]
  reg [21:0] _T_3632; // @[Reg.scala 27:20]
  reg [21:0] _T_3571; // @[Reg.scala 27:20]
  reg [21:0] _T_3510; // @[Reg.scala 27:20]
  reg [21:0] _T_3449; // @[Reg.scala 27:20]
  reg [21:0] _T_3388; // @[Reg.scala 27:20]
  reg [21:0] _T_3327; // @[Reg.scala 27:20]
  reg [21:0] _T_3266; // @[Reg.scala 27:20]
  reg [21:0] _T_3205; // @[Reg.scala 27:20]
  reg [21:0] _T_3144; // @[Reg.scala 27:20]
  reg [21:0] _T_3083; // @[Reg.scala 27:20]
  reg [21:0] _T_3022; // @[Reg.scala 27:20]
  reg [21:0] _T_2961; // @[Reg.scala 27:20]
  reg [21:0] _T_2900; // @[Reg.scala 27:20]
  reg [21:0] _T_2839; // @[Reg.scala 27:20]
  reg [21:0] _T_2778; // @[Reg.scala 27:20]
  reg [21:0] _T_2717; // @[Reg.scala 27:20]
  reg [21:0] _T_2656; // @[Reg.scala 27:20]
  reg [21:0] _T_2595; // @[Reg.scala 27:20]
  reg [21:0] _T_2534; // @[Reg.scala 27:20]
  reg [21:0] _T_2473; // @[Reg.scala 27:20]
  reg [21:0] _T_2412; // @[Reg.scala 27:20]
  reg [21:0] _T_2351; // @[Reg.scala 27:20]
  reg [21:0] _T_2290; // @[Reg.scala 27:20]
  reg [21:0] _T_2229; // @[Reg.scala 27:20]
  reg [21:0] _T_2168; // @[Reg.scala 27:20]
  reg [21:0] _T_2107; // @[Reg.scala 27:20]
  reg [21:0] _T_2046; // @[Reg.scala 27:20]
  reg [21:0] _T_1985; // @[Reg.scala 27:20]
  reg [21:0] _T_1924; // @[Reg.scala 27:20]
  reg [21:0] _T_1863; // @[Reg.scala 27:20]
  reg [21:0] _T_1802; // @[Reg.scala 27:20]
  reg [21:0] _T_1741; // @[Reg.scala 27:20]
  reg [21:0] _T_1680; // @[Reg.scala 27:20]
  reg [21:0] _T_1619; // @[Reg.scala 27:20]
  reg [21:0] _T_1558; // @[Reg.scala 27:20]
  reg [21:0] _T_1497; // @[Reg.scala 27:20]
  reg [21:0] _T_1436; // @[Reg.scala 27:20]
  reg [21:0] _T_1375; // @[Reg.scala 27:20]
  reg [21:0] _T_1314; // @[Reg.scala 27:20]
  reg [21:0] _T_1253; // @[Reg.scala 27:20]
  reg [21:0] _T_1192; // @[Reg.scala 27:20]
  reg [21:0] _T_1131; // @[Reg.scala 27:20]
  reg [21:0] _T_1070; // @[Reg.scala 27:20]
  reg [21:0] _T_1009; // @[Reg.scala 27:20]
  reg [21:0] _T_948; // @[Reg.scala 27:20]
  reg [21:0] _T_887; // @[Reg.scala 27:20]
  reg [21:0] _T_826; // @[Reg.scala 27:20]
  reg [21:0] _T_765; // @[Reg.scala 27:20]
  reg [21:0] _T_704; // @[Reg.scala 27:20]
  reg [21:0] _T_643; // @[Reg.scala 27:20]
  reg [21:0] _T_582; // @[Reg.scala 27:20]
  reg [21:0] _T_521; // @[Reg.scala 27:20]
  reg [21:0] _T_460; // @[Reg.scala 27:20]
  wire [21:0] _T_32_1 = _T_157 ? _T_521 : _T_460; // @[Mux.scala 80:57]
  wire [21:0] _T_34_1 = _T_159 ? _T_582 : _T_32_1; // @[Mux.scala 80:57]
  wire [21:0] _T_36_1 = _T_161 ? _T_643 : _T_34_1; // @[Mux.scala 80:57]
  wire [21:0] _T_38_1 = _T_163 ? _T_704 : _T_36_1; // @[Mux.scala 80:57]
  wire [21:0] _T_40_1 = _T_165 ? _T_765 : _T_38_1; // @[Mux.scala 80:57]
  wire [21:0] _T_42_1 = _T_167 ? _T_826 : _T_40_1; // @[Mux.scala 80:57]
  wire [21:0] _T_44_1 = _T_169 ? _T_887 : _T_42_1; // @[Mux.scala 80:57]
  wire [21:0] _T_46_1 = _T_171 ? _T_948 : _T_44_1; // @[Mux.scala 80:57]
  wire [21:0] _T_48_1 = _T_173 ? _T_1009 : _T_46_1; // @[Mux.scala 80:57]
  wire [21:0] _T_50_1 = _T_175 ? _T_1070 : _T_48_1; // @[Mux.scala 80:57]
  wire [21:0] _T_52_1 = _T_177 ? _T_1131 : _T_50_1; // @[Mux.scala 80:57]
  wire [21:0] _T_54_1 = _T_179 ? _T_1192 : _T_52_1; // @[Mux.scala 80:57]
  wire [21:0] _T_56_1 = _T_181 ? _T_1253 : _T_54_1; // @[Mux.scala 80:57]
  wire [21:0] _T_58_1 = _T_183 ? _T_1314 : _T_56_1; // @[Mux.scala 80:57]
  wire [21:0] _T_60_1 = _T_185 ? _T_1375 : _T_58_1; // @[Mux.scala 80:57]
  wire [21:0] _T_62_1 = _T_187 ? _T_1436 : _T_60_1; // @[Mux.scala 80:57]
  wire [21:0] _T_64_1 = _T_189 ? _T_1497 : _T_62_1; // @[Mux.scala 80:57]
  wire [21:0] _T_66_1 = _T_191 ? _T_1558 : _T_64_1; // @[Mux.scala 80:57]
  wire [21:0] _T_68_1 = _T_193 ? _T_1619 : _T_66_1; // @[Mux.scala 80:57]
  wire [21:0] _T_70_1 = _T_195 ? _T_1680 : _T_68_1; // @[Mux.scala 80:57]
  wire [21:0] _T_72_1 = _T_197 ? _T_1741 : _T_70_1; // @[Mux.scala 80:57]
  wire [21:0] _T_74_1 = _T_199 ? _T_1802 : _T_72_1; // @[Mux.scala 80:57]
  wire [21:0] _T_76_1 = _T_201 ? _T_1863 : _T_74_1; // @[Mux.scala 80:57]
  wire [21:0] _T_78_1 = _T_203 ? _T_1924 : _T_76_1; // @[Mux.scala 80:57]
  wire [21:0] _T_80_1 = _T_205 ? _T_1985 : _T_78_1; // @[Mux.scala 80:57]
  wire [21:0] _T_82_1 = _T_207 ? _T_2046 : _T_80_1; // @[Mux.scala 80:57]
  wire [21:0] _T_84_1 = _T_209 ? _T_2107 : _T_82_1; // @[Mux.scala 80:57]
  wire [21:0] _T_86_1 = _T_211 ? _T_2168 : _T_84_1; // @[Mux.scala 80:57]
  wire [21:0] _T_88_1 = _T_213 ? _T_2229 : _T_86_1; // @[Mux.scala 80:57]
  wire [21:0] _T_90_1 = _T_215 ? _T_2290 : _T_88_1; // @[Mux.scala 80:57]
  wire [21:0] _T_92_1 = _T_217 ? _T_2351 : _T_90_1; // @[Mux.scala 80:57]
  wire [21:0] _T_94_1 = _T_219 ? _T_2412 : _T_92_1; // @[Mux.scala 80:57]
  wire [21:0] _T_96_1 = _T_221 ? _T_2473 : _T_94_1; // @[Mux.scala 80:57]
  wire [21:0] _T_98_1 = _T_223 ? _T_2534 : _T_96_1; // @[Mux.scala 80:57]
  wire [21:0] _T_100_1 = _T_225 ? _T_2595 : _T_98_1; // @[Mux.scala 80:57]
  wire [21:0] _T_102_1 = _T_227 ? _T_2656 : _T_100_1; // @[Mux.scala 80:57]
  wire [21:0] _T_104_1 = _T_229 ? _T_2717 : _T_102_1; // @[Mux.scala 80:57]
  wire [21:0] _T_106_1 = _T_231 ? _T_2778 : _T_104_1; // @[Mux.scala 80:57]
  wire [21:0] _T_108_1 = _T_233 ? _T_2839 : _T_106_1; // @[Mux.scala 80:57]
  wire [21:0] _T_110_1 = _T_235 ? _T_2900 : _T_108_1; // @[Mux.scala 80:57]
  wire [21:0] _T_112_1 = _T_237 ? _T_2961 : _T_110_1; // @[Mux.scala 80:57]
  wire [21:0] _T_114_1 = _T_239 ? _T_3022 : _T_112_1; // @[Mux.scala 80:57]
  wire [21:0] _T_116_1 = _T_241 ? _T_3083 : _T_114_1; // @[Mux.scala 80:57]
  wire [21:0] _T_118_1 = _T_243 ? _T_3144 : _T_116_1; // @[Mux.scala 80:57]
  wire [21:0] _T_120_1 = _T_245 ? _T_3205 : _T_118_1; // @[Mux.scala 80:57]
  wire [21:0] _T_122_1 = _T_247 ? _T_3266 : _T_120_1; // @[Mux.scala 80:57]
  wire [21:0] _T_124_1 = _T_249 ? _T_3327 : _T_122_1; // @[Mux.scala 80:57]
  wire [21:0] _T_126_1 = _T_251 ? _T_3388 : _T_124_1; // @[Mux.scala 80:57]
  wire [21:0] _T_128_1 = _T_253 ? _T_3449 : _T_126_1; // @[Mux.scala 80:57]
  wire [21:0] _T_130_1 = _T_255 ? _T_3510 : _T_128_1; // @[Mux.scala 80:57]
  wire [21:0] _T_132_1 = _T_257 ? _T_3571 : _T_130_1; // @[Mux.scala 80:57]
  wire [21:0] _T_134_1 = _T_259 ? _T_3632 : _T_132_1; // @[Mux.scala 80:57]
  wire [21:0] _T_136_1 = _T_261 ? _T_3693 : _T_134_1; // @[Mux.scala 80:57]
  wire [21:0] _T_138_1 = _T_263 ? _T_3754 : _T_136_1; // @[Mux.scala 80:57]
  wire [21:0] _T_140_1 = _T_265 ? _T_3815 : _T_138_1; // @[Mux.scala 80:57]
  wire [21:0] _T_142_1 = _T_267 ? _T_3876 : _T_140_1; // @[Mux.scala 80:57]
  wire [21:0] _T_144_1 = _T_269 ? _T_3937 : _T_142_1; // @[Mux.scala 80:57]
  wire [21:0] _T_146_1 = _T_271 ? _T_3998 : _T_144_1; // @[Mux.scala 80:57]
  wire [21:0] _T_148_1 = _T_273 ? _T_4059 : _T_146_1; // @[Mux.scala 80:57]
  wire [21:0] _T_150_1 = _T_275 ? _T_4120 : _T_148_1; // @[Mux.scala 80:57]
  wire [21:0] _T_152_1 = _T_277 ? _T_4181 : _T_150_1; // @[Mux.scala 80:57]
  wire [21:0] _T_154_1 = _T_279 ? _T_4242 : _T_152_1; // @[Mux.scala 80:57]
  wire [21:0] _T_156_1 = _T_281 ? _T_4303 : _T_154_1; // @[Mux.scala 80:57]
  wire  _T_285 = _T_156_1 == io_cacheIn_addr[31:10]; // @[Cache.scala 772:78]
  wire  _T_286 = _T_282_1 & _T_285; // @[Cache.scala 772:62]
  wire  _T_292 = _T_284 | _T_286; // @[Cache.scala 773:51]
  reg  _T_4325; // @[Reg.scala 27:20]
  reg  _T_4264; // @[Reg.scala 27:20]
  reg  _T_4203; // @[Reg.scala 27:20]
  reg  _T_4142; // @[Reg.scala 27:20]
  reg  _T_4081; // @[Reg.scala 27:20]
  reg  _T_4020; // @[Reg.scala 27:20]
  reg  _T_3959; // @[Reg.scala 27:20]
  reg  _T_3898; // @[Reg.scala 27:20]
  reg  _T_3837; // @[Reg.scala 27:20]
  reg  _T_3776; // @[Reg.scala 27:20]
  reg  _T_3715; // @[Reg.scala 27:20]
  reg  _T_3654; // @[Reg.scala 27:20]
  reg  _T_3593; // @[Reg.scala 27:20]
  reg  _T_3532; // @[Reg.scala 27:20]
  reg  _T_3471; // @[Reg.scala 27:20]
  reg  _T_3410; // @[Reg.scala 27:20]
  reg  _T_3349; // @[Reg.scala 27:20]
  reg  _T_3288; // @[Reg.scala 27:20]
  reg  _T_3227; // @[Reg.scala 27:20]
  reg  _T_3166; // @[Reg.scala 27:20]
  reg  _T_3105; // @[Reg.scala 27:20]
  reg  _T_3044; // @[Reg.scala 27:20]
  reg  _T_2983; // @[Reg.scala 27:20]
  reg  _T_2922; // @[Reg.scala 27:20]
  reg  _T_2861; // @[Reg.scala 27:20]
  reg  _T_2800; // @[Reg.scala 27:20]
  reg  _T_2739; // @[Reg.scala 27:20]
  reg  _T_2678; // @[Reg.scala 27:20]
  reg  _T_2617; // @[Reg.scala 27:20]
  reg  _T_2556; // @[Reg.scala 27:20]
  reg  _T_2495; // @[Reg.scala 27:20]
  reg  _T_2434; // @[Reg.scala 27:20]
  reg  _T_2373; // @[Reg.scala 27:20]
  reg  _T_2312; // @[Reg.scala 27:20]
  reg  _T_2251; // @[Reg.scala 27:20]
  reg  _T_2190; // @[Reg.scala 27:20]
  reg  _T_2129; // @[Reg.scala 27:20]
  reg  _T_2068; // @[Reg.scala 27:20]
  reg  _T_2007; // @[Reg.scala 27:20]
  reg  _T_1946; // @[Reg.scala 27:20]
  reg  _T_1885; // @[Reg.scala 27:20]
  reg  _T_1824; // @[Reg.scala 27:20]
  reg  _T_1763; // @[Reg.scala 27:20]
  reg  _T_1702; // @[Reg.scala 27:20]
  reg  _T_1641; // @[Reg.scala 27:20]
  reg  _T_1580; // @[Reg.scala 27:20]
  reg  _T_1519; // @[Reg.scala 27:20]
  reg  _T_1458; // @[Reg.scala 27:20]
  reg  _T_1397; // @[Reg.scala 27:20]
  reg  _T_1336; // @[Reg.scala 27:20]
  reg  _T_1275; // @[Reg.scala 27:20]
  reg  _T_1214; // @[Reg.scala 27:20]
  reg  _T_1153; // @[Reg.scala 27:20]
  reg  _T_1092; // @[Reg.scala 27:20]
  reg  _T_1031; // @[Reg.scala 27:20]
  reg  _T_970; // @[Reg.scala 27:20]
  reg  _T_909; // @[Reg.scala 27:20]
  reg  _T_848; // @[Reg.scala 27:20]
  reg  _T_787; // @[Reg.scala 27:20]
  reg  _T_726; // @[Reg.scala 27:20]
  reg  _T_665; // @[Reg.scala 27:20]
  reg  _T_604; // @[Reg.scala 27:20]
  reg  _T_543; // @[Reg.scala 27:20]
  reg  _T_482; // @[Reg.scala 27:20]
  wire  _T_158_2 = _T_157 ? _T_543 : _T_482; // @[Mux.scala 80:57]
  wire  _T_160_2 = _T_159 ? _T_604 : _T_158_2; // @[Mux.scala 80:57]
  wire  _T_162_2 = _T_161 ? _T_665 : _T_160_2; // @[Mux.scala 80:57]
  wire  _T_164_2 = _T_163 ? _T_726 : _T_162_2; // @[Mux.scala 80:57]
  wire  _T_166_2 = _T_165 ? _T_787 : _T_164_2; // @[Mux.scala 80:57]
  wire  _T_168_2 = _T_167 ? _T_848 : _T_166_2; // @[Mux.scala 80:57]
  wire  _T_170_2 = _T_169 ? _T_909 : _T_168_2; // @[Mux.scala 80:57]
  wire  _T_172_2 = _T_171 ? _T_970 : _T_170_2; // @[Mux.scala 80:57]
  wire  _T_174_2 = _T_173 ? _T_1031 : _T_172_2; // @[Mux.scala 80:57]
  wire  _T_176_2 = _T_175 ? _T_1092 : _T_174_2; // @[Mux.scala 80:57]
  wire  _T_178_2 = _T_177 ? _T_1153 : _T_176_2; // @[Mux.scala 80:57]
  wire  _T_180_2 = _T_179 ? _T_1214 : _T_178_2; // @[Mux.scala 80:57]
  wire  _T_182_2 = _T_181 ? _T_1275 : _T_180_2; // @[Mux.scala 80:57]
  wire  _T_184_2 = _T_183 ? _T_1336 : _T_182_2; // @[Mux.scala 80:57]
  wire  _T_186_2 = _T_185 ? _T_1397 : _T_184_2; // @[Mux.scala 80:57]
  wire  _T_188_2 = _T_187 ? _T_1458 : _T_186_2; // @[Mux.scala 80:57]
  wire  _T_190_2 = _T_189 ? _T_1519 : _T_188_2; // @[Mux.scala 80:57]
  wire  _T_192_2 = _T_191 ? _T_1580 : _T_190_2; // @[Mux.scala 80:57]
  wire  _T_194_2 = _T_193 ? _T_1641 : _T_192_2; // @[Mux.scala 80:57]
  wire  _T_196_2 = _T_195 ? _T_1702 : _T_194_2; // @[Mux.scala 80:57]
  wire  _T_198_2 = _T_197 ? _T_1763 : _T_196_2; // @[Mux.scala 80:57]
  wire  _T_200_2 = _T_199 ? _T_1824 : _T_198_2; // @[Mux.scala 80:57]
  wire  _T_202_2 = _T_201 ? _T_1885 : _T_200_2; // @[Mux.scala 80:57]
  wire  _T_204_2 = _T_203 ? _T_1946 : _T_202_2; // @[Mux.scala 80:57]
  wire  _T_206_2 = _T_205 ? _T_2007 : _T_204_2; // @[Mux.scala 80:57]
  wire  _T_208_2 = _T_207 ? _T_2068 : _T_206_2; // @[Mux.scala 80:57]
  wire  _T_210_2 = _T_209 ? _T_2129 : _T_208_2; // @[Mux.scala 80:57]
  wire  _T_212_2 = _T_211 ? _T_2190 : _T_210_2; // @[Mux.scala 80:57]
  wire  _T_214_2 = _T_213 ? _T_2251 : _T_212_2; // @[Mux.scala 80:57]
  wire  _T_216_2 = _T_215 ? _T_2312 : _T_214_2; // @[Mux.scala 80:57]
  wire  _T_218_2 = _T_217 ? _T_2373 : _T_216_2; // @[Mux.scala 80:57]
  wire  _T_220_2 = _T_219 ? _T_2434 : _T_218_2; // @[Mux.scala 80:57]
  wire  _T_222_2 = _T_221 ? _T_2495 : _T_220_2; // @[Mux.scala 80:57]
  wire  _T_224_2 = _T_223 ? _T_2556 : _T_222_2; // @[Mux.scala 80:57]
  wire  _T_226_2 = _T_225 ? _T_2617 : _T_224_2; // @[Mux.scala 80:57]
  wire  _T_228_2 = _T_227 ? _T_2678 : _T_226_2; // @[Mux.scala 80:57]
  wire  _T_230_2 = _T_229 ? _T_2739 : _T_228_2; // @[Mux.scala 80:57]
  wire  _T_232_2 = _T_231 ? _T_2800 : _T_230_2; // @[Mux.scala 80:57]
  wire  _T_234_2 = _T_233 ? _T_2861 : _T_232_2; // @[Mux.scala 80:57]
  wire  _T_236_2 = _T_235 ? _T_2922 : _T_234_2; // @[Mux.scala 80:57]
  wire  _T_238_2 = _T_237 ? _T_2983 : _T_236_2; // @[Mux.scala 80:57]
  wire  _T_240_2 = _T_239 ? _T_3044 : _T_238_2; // @[Mux.scala 80:57]
  wire  _T_242_2 = _T_241 ? _T_3105 : _T_240_2; // @[Mux.scala 80:57]
  wire  _T_244_2 = _T_243 ? _T_3166 : _T_242_2; // @[Mux.scala 80:57]
  wire  _T_246_2 = _T_245 ? _T_3227 : _T_244_2; // @[Mux.scala 80:57]
  wire  _T_248_2 = _T_247 ? _T_3288 : _T_246_2; // @[Mux.scala 80:57]
  wire  _T_250_2 = _T_249 ? _T_3349 : _T_248_2; // @[Mux.scala 80:57]
  wire  _T_252_2 = _T_251 ? _T_3410 : _T_250_2; // @[Mux.scala 80:57]
  wire  _T_254_2 = _T_253 ? _T_3471 : _T_252_2; // @[Mux.scala 80:57]
  wire  _T_256_2 = _T_255 ? _T_3532 : _T_254_2; // @[Mux.scala 80:57]
  wire  _T_258_2 = _T_257 ? _T_3593 : _T_256_2; // @[Mux.scala 80:57]
  wire  _T_260_2 = _T_259 ? _T_3654 : _T_258_2; // @[Mux.scala 80:57]
  wire  _T_262_2 = _T_261 ? _T_3715 : _T_260_2; // @[Mux.scala 80:57]
  wire  _T_264_2 = _T_263 ? _T_3776 : _T_262_2; // @[Mux.scala 80:57]
  wire  _T_266_2 = _T_265 ? _T_3837 : _T_264_2; // @[Mux.scala 80:57]
  wire  _T_268_2 = _T_267 ? _T_3898 : _T_266_2; // @[Mux.scala 80:57]
  wire  _T_270_2 = _T_269 ? _T_3959 : _T_268_2; // @[Mux.scala 80:57]
  wire  _T_272_2 = _T_271 ? _T_4020 : _T_270_2; // @[Mux.scala 80:57]
  wire  _T_274_2 = _T_273 ? _T_4081 : _T_272_2; // @[Mux.scala 80:57]
  wire  _T_276_2 = _T_275 ? _T_4142 : _T_274_2; // @[Mux.scala 80:57]
  wire  _T_278_2 = _T_277 ? _T_4203 : _T_276_2; // @[Mux.scala 80:57]
  wire  _T_280_2 = _T_279 ? _T_4264 : _T_278_2; // @[Mux.scala 80:57]
  wire  _T_282_2 = _T_281 ? _T_4325 : _T_280_2; // @[Mux.scala 80:57]
  reg [21:0] _T_4317; // @[Reg.scala 27:20]
  reg [21:0] _T_4256; // @[Reg.scala 27:20]
  reg [21:0] _T_4195; // @[Reg.scala 27:20]
  reg [21:0] _T_4134; // @[Reg.scala 27:20]
  reg [21:0] _T_4073; // @[Reg.scala 27:20]
  reg [21:0] _T_4012; // @[Reg.scala 27:20]
  reg [21:0] _T_3951; // @[Reg.scala 27:20]
  reg [21:0] _T_3890; // @[Reg.scala 27:20]
  reg [21:0] _T_3829; // @[Reg.scala 27:20]
  reg [21:0] _T_3768; // @[Reg.scala 27:20]
  reg [21:0] _T_3707; // @[Reg.scala 27:20]
  reg [21:0] _T_3646; // @[Reg.scala 27:20]
  reg [21:0] _T_3585; // @[Reg.scala 27:20]
  reg [21:0] _T_3524; // @[Reg.scala 27:20]
  reg [21:0] _T_3463; // @[Reg.scala 27:20]
  reg [21:0] _T_3402; // @[Reg.scala 27:20]
  reg [21:0] _T_3341; // @[Reg.scala 27:20]
  reg [21:0] _T_3280; // @[Reg.scala 27:20]
  reg [21:0] _T_3219; // @[Reg.scala 27:20]
  reg [21:0] _T_3158; // @[Reg.scala 27:20]
  reg [21:0] _T_3097; // @[Reg.scala 27:20]
  reg [21:0] _T_3036; // @[Reg.scala 27:20]
  reg [21:0] _T_2975; // @[Reg.scala 27:20]
  reg [21:0] _T_2914; // @[Reg.scala 27:20]
  reg [21:0] _T_2853; // @[Reg.scala 27:20]
  reg [21:0] _T_2792; // @[Reg.scala 27:20]
  reg [21:0] _T_2731; // @[Reg.scala 27:20]
  reg [21:0] _T_2670; // @[Reg.scala 27:20]
  reg [21:0] _T_2609; // @[Reg.scala 27:20]
  reg [21:0] _T_2548; // @[Reg.scala 27:20]
  reg [21:0] _T_2487; // @[Reg.scala 27:20]
  reg [21:0] _T_2426; // @[Reg.scala 27:20]
  reg [21:0] _T_2365; // @[Reg.scala 27:20]
  reg [21:0] _T_2304; // @[Reg.scala 27:20]
  reg [21:0] _T_2243; // @[Reg.scala 27:20]
  reg [21:0] _T_2182; // @[Reg.scala 27:20]
  reg [21:0] _T_2121; // @[Reg.scala 27:20]
  reg [21:0] _T_2060; // @[Reg.scala 27:20]
  reg [21:0] _T_1999; // @[Reg.scala 27:20]
  reg [21:0] _T_1938; // @[Reg.scala 27:20]
  reg [21:0] _T_1877; // @[Reg.scala 27:20]
  reg [21:0] _T_1816; // @[Reg.scala 27:20]
  reg [21:0] _T_1755; // @[Reg.scala 27:20]
  reg [21:0] _T_1694; // @[Reg.scala 27:20]
  reg [21:0] _T_1633; // @[Reg.scala 27:20]
  reg [21:0] _T_1572; // @[Reg.scala 27:20]
  reg [21:0] _T_1511; // @[Reg.scala 27:20]
  reg [21:0] _T_1450; // @[Reg.scala 27:20]
  reg [21:0] _T_1389; // @[Reg.scala 27:20]
  reg [21:0] _T_1328; // @[Reg.scala 27:20]
  reg [21:0] _T_1267; // @[Reg.scala 27:20]
  reg [21:0] _T_1206; // @[Reg.scala 27:20]
  reg [21:0] _T_1145; // @[Reg.scala 27:20]
  reg [21:0] _T_1084; // @[Reg.scala 27:20]
  reg [21:0] _T_1023; // @[Reg.scala 27:20]
  reg [21:0] _T_962; // @[Reg.scala 27:20]
  reg [21:0] _T_901; // @[Reg.scala 27:20]
  reg [21:0] _T_840; // @[Reg.scala 27:20]
  reg [21:0] _T_779; // @[Reg.scala 27:20]
  reg [21:0] _T_718; // @[Reg.scala 27:20]
  reg [21:0] _T_657; // @[Reg.scala 27:20]
  reg [21:0] _T_596; // @[Reg.scala 27:20]
  reg [21:0] _T_535; // @[Reg.scala 27:20]
  reg [21:0] _T_474; // @[Reg.scala 27:20]
  wire [21:0] _T_32_2 = _T_157 ? _T_535 : _T_474; // @[Mux.scala 80:57]
  wire [21:0] _T_34_2 = _T_159 ? _T_596 : _T_32_2; // @[Mux.scala 80:57]
  wire [21:0] _T_36_2 = _T_161 ? _T_657 : _T_34_2; // @[Mux.scala 80:57]
  wire [21:0] _T_38_2 = _T_163 ? _T_718 : _T_36_2; // @[Mux.scala 80:57]
  wire [21:0] _T_40_2 = _T_165 ? _T_779 : _T_38_2; // @[Mux.scala 80:57]
  wire [21:0] _T_42_2 = _T_167 ? _T_840 : _T_40_2; // @[Mux.scala 80:57]
  wire [21:0] _T_44_2 = _T_169 ? _T_901 : _T_42_2; // @[Mux.scala 80:57]
  wire [21:0] _T_46_2 = _T_171 ? _T_962 : _T_44_2; // @[Mux.scala 80:57]
  wire [21:0] _T_48_2 = _T_173 ? _T_1023 : _T_46_2; // @[Mux.scala 80:57]
  wire [21:0] _T_50_2 = _T_175 ? _T_1084 : _T_48_2; // @[Mux.scala 80:57]
  wire [21:0] _T_52_2 = _T_177 ? _T_1145 : _T_50_2; // @[Mux.scala 80:57]
  wire [21:0] _T_54_2 = _T_179 ? _T_1206 : _T_52_2; // @[Mux.scala 80:57]
  wire [21:0] _T_56_2 = _T_181 ? _T_1267 : _T_54_2; // @[Mux.scala 80:57]
  wire [21:0] _T_58_2 = _T_183 ? _T_1328 : _T_56_2; // @[Mux.scala 80:57]
  wire [21:0] _T_60_2 = _T_185 ? _T_1389 : _T_58_2; // @[Mux.scala 80:57]
  wire [21:0] _T_62_2 = _T_187 ? _T_1450 : _T_60_2; // @[Mux.scala 80:57]
  wire [21:0] _T_64_2 = _T_189 ? _T_1511 : _T_62_2; // @[Mux.scala 80:57]
  wire [21:0] _T_66_2 = _T_191 ? _T_1572 : _T_64_2; // @[Mux.scala 80:57]
  wire [21:0] _T_68_2 = _T_193 ? _T_1633 : _T_66_2; // @[Mux.scala 80:57]
  wire [21:0] _T_70_2 = _T_195 ? _T_1694 : _T_68_2; // @[Mux.scala 80:57]
  wire [21:0] _T_72_2 = _T_197 ? _T_1755 : _T_70_2; // @[Mux.scala 80:57]
  wire [21:0] _T_74_2 = _T_199 ? _T_1816 : _T_72_2; // @[Mux.scala 80:57]
  wire [21:0] _T_76_2 = _T_201 ? _T_1877 : _T_74_2; // @[Mux.scala 80:57]
  wire [21:0] _T_78_2 = _T_203 ? _T_1938 : _T_76_2; // @[Mux.scala 80:57]
  wire [21:0] _T_80_2 = _T_205 ? _T_1999 : _T_78_2; // @[Mux.scala 80:57]
  wire [21:0] _T_82_2 = _T_207 ? _T_2060 : _T_80_2; // @[Mux.scala 80:57]
  wire [21:0] _T_84_2 = _T_209 ? _T_2121 : _T_82_2; // @[Mux.scala 80:57]
  wire [21:0] _T_86_2 = _T_211 ? _T_2182 : _T_84_2; // @[Mux.scala 80:57]
  wire [21:0] _T_88_2 = _T_213 ? _T_2243 : _T_86_2; // @[Mux.scala 80:57]
  wire [21:0] _T_90_2 = _T_215 ? _T_2304 : _T_88_2; // @[Mux.scala 80:57]
  wire [21:0] _T_92_2 = _T_217 ? _T_2365 : _T_90_2; // @[Mux.scala 80:57]
  wire [21:0] _T_94_2 = _T_219 ? _T_2426 : _T_92_2; // @[Mux.scala 80:57]
  wire [21:0] _T_96_2 = _T_221 ? _T_2487 : _T_94_2; // @[Mux.scala 80:57]
  wire [21:0] _T_98_2 = _T_223 ? _T_2548 : _T_96_2; // @[Mux.scala 80:57]
  wire [21:0] _T_100_2 = _T_225 ? _T_2609 : _T_98_2; // @[Mux.scala 80:57]
  wire [21:0] _T_102_2 = _T_227 ? _T_2670 : _T_100_2; // @[Mux.scala 80:57]
  wire [21:0] _T_104_2 = _T_229 ? _T_2731 : _T_102_2; // @[Mux.scala 80:57]
  wire [21:0] _T_106_2 = _T_231 ? _T_2792 : _T_104_2; // @[Mux.scala 80:57]
  wire [21:0] _T_108_2 = _T_233 ? _T_2853 : _T_106_2; // @[Mux.scala 80:57]
  wire [21:0] _T_110_2 = _T_235 ? _T_2914 : _T_108_2; // @[Mux.scala 80:57]
  wire [21:0] _T_112_2 = _T_237 ? _T_2975 : _T_110_2; // @[Mux.scala 80:57]
  wire [21:0] _T_114_2 = _T_239 ? _T_3036 : _T_112_2; // @[Mux.scala 80:57]
  wire [21:0] _T_116_2 = _T_241 ? _T_3097 : _T_114_2; // @[Mux.scala 80:57]
  wire [21:0] _T_118_2 = _T_243 ? _T_3158 : _T_116_2; // @[Mux.scala 80:57]
  wire [21:0] _T_120_2 = _T_245 ? _T_3219 : _T_118_2; // @[Mux.scala 80:57]
  wire [21:0] _T_122_2 = _T_247 ? _T_3280 : _T_120_2; // @[Mux.scala 80:57]
  wire [21:0] _T_124_2 = _T_249 ? _T_3341 : _T_122_2; // @[Mux.scala 80:57]
  wire [21:0] _T_126_2 = _T_251 ? _T_3402 : _T_124_2; // @[Mux.scala 80:57]
  wire [21:0] _T_128_2 = _T_253 ? _T_3463 : _T_126_2; // @[Mux.scala 80:57]
  wire [21:0] _T_130_2 = _T_255 ? _T_3524 : _T_128_2; // @[Mux.scala 80:57]
  wire [21:0] _T_132_2 = _T_257 ? _T_3585 : _T_130_2; // @[Mux.scala 80:57]
  wire [21:0] _T_134_2 = _T_259 ? _T_3646 : _T_132_2; // @[Mux.scala 80:57]
  wire [21:0] _T_136_2 = _T_261 ? _T_3707 : _T_134_2; // @[Mux.scala 80:57]
  wire [21:0] _T_138_2 = _T_263 ? _T_3768 : _T_136_2; // @[Mux.scala 80:57]
  wire [21:0] _T_140_2 = _T_265 ? _T_3829 : _T_138_2; // @[Mux.scala 80:57]
  wire [21:0] _T_142_2 = _T_267 ? _T_3890 : _T_140_2; // @[Mux.scala 80:57]
  wire [21:0] _T_144_2 = _T_269 ? _T_3951 : _T_142_2; // @[Mux.scala 80:57]
  wire [21:0] _T_146_2 = _T_271 ? _T_4012 : _T_144_2; // @[Mux.scala 80:57]
  wire [21:0] _T_148_2 = _T_273 ? _T_4073 : _T_146_2; // @[Mux.scala 80:57]
  wire [21:0] _T_150_2 = _T_275 ? _T_4134 : _T_148_2; // @[Mux.scala 80:57]
  wire [21:0] _T_152_2 = _T_277 ? _T_4195 : _T_150_2; // @[Mux.scala 80:57]
  wire [21:0] _T_154_2 = _T_279 ? _T_4256 : _T_152_2; // @[Mux.scala 80:57]
  wire [21:0] _T_156_2 = _T_281 ? _T_4317 : _T_154_2; // @[Mux.scala 80:57]
  wire  _T_287 = _T_156_2 == io_cacheIn_addr[31:10]; // @[Cache.scala 772:78]
  wire  _T_288 = _T_282_2 & _T_287; // @[Cache.scala 772:62]
  wire  _T_293 = _T_292 | _T_288; // @[Cache.scala 773:51]
  reg  _T_4339; // @[Reg.scala 27:20]
  reg  _T_4278; // @[Reg.scala 27:20]
  reg  _T_4217; // @[Reg.scala 27:20]
  reg  _T_4156; // @[Reg.scala 27:20]
  reg  _T_4095; // @[Reg.scala 27:20]
  reg  _T_4034; // @[Reg.scala 27:20]
  reg  _T_3973; // @[Reg.scala 27:20]
  reg  _T_3912; // @[Reg.scala 27:20]
  reg  _T_3851; // @[Reg.scala 27:20]
  reg  _T_3790; // @[Reg.scala 27:20]
  reg  _T_3729; // @[Reg.scala 27:20]
  reg  _T_3668; // @[Reg.scala 27:20]
  reg  _T_3607; // @[Reg.scala 27:20]
  reg  _T_3546; // @[Reg.scala 27:20]
  reg  _T_3485; // @[Reg.scala 27:20]
  reg  _T_3424; // @[Reg.scala 27:20]
  reg  _T_3363; // @[Reg.scala 27:20]
  reg  _T_3302; // @[Reg.scala 27:20]
  reg  _T_3241; // @[Reg.scala 27:20]
  reg  _T_3180; // @[Reg.scala 27:20]
  reg  _T_3119; // @[Reg.scala 27:20]
  reg  _T_3058; // @[Reg.scala 27:20]
  reg  _T_2997; // @[Reg.scala 27:20]
  reg  _T_2936; // @[Reg.scala 27:20]
  reg  _T_2875; // @[Reg.scala 27:20]
  reg  _T_2814; // @[Reg.scala 27:20]
  reg  _T_2753; // @[Reg.scala 27:20]
  reg  _T_2692; // @[Reg.scala 27:20]
  reg  _T_2631; // @[Reg.scala 27:20]
  reg  _T_2570; // @[Reg.scala 27:20]
  reg  _T_2509; // @[Reg.scala 27:20]
  reg  _T_2448; // @[Reg.scala 27:20]
  reg  _T_2387; // @[Reg.scala 27:20]
  reg  _T_2326; // @[Reg.scala 27:20]
  reg  _T_2265; // @[Reg.scala 27:20]
  reg  _T_2204; // @[Reg.scala 27:20]
  reg  _T_2143; // @[Reg.scala 27:20]
  reg  _T_2082; // @[Reg.scala 27:20]
  reg  _T_2021; // @[Reg.scala 27:20]
  reg  _T_1960; // @[Reg.scala 27:20]
  reg  _T_1899; // @[Reg.scala 27:20]
  reg  _T_1838; // @[Reg.scala 27:20]
  reg  _T_1777; // @[Reg.scala 27:20]
  reg  _T_1716; // @[Reg.scala 27:20]
  reg  _T_1655; // @[Reg.scala 27:20]
  reg  _T_1594; // @[Reg.scala 27:20]
  reg  _T_1533; // @[Reg.scala 27:20]
  reg  _T_1472; // @[Reg.scala 27:20]
  reg  _T_1411; // @[Reg.scala 27:20]
  reg  _T_1350; // @[Reg.scala 27:20]
  reg  _T_1289; // @[Reg.scala 27:20]
  reg  _T_1228; // @[Reg.scala 27:20]
  reg  _T_1167; // @[Reg.scala 27:20]
  reg  _T_1106; // @[Reg.scala 27:20]
  reg  _T_1045; // @[Reg.scala 27:20]
  reg  _T_984; // @[Reg.scala 27:20]
  reg  _T_923; // @[Reg.scala 27:20]
  reg  _T_862; // @[Reg.scala 27:20]
  reg  _T_801; // @[Reg.scala 27:20]
  reg  _T_740; // @[Reg.scala 27:20]
  reg  _T_679; // @[Reg.scala 27:20]
  reg  _T_618; // @[Reg.scala 27:20]
  reg  _T_557; // @[Reg.scala 27:20]
  reg  _T_496; // @[Reg.scala 27:20]
  wire  _T_158_3 = _T_157 ? _T_557 : _T_496; // @[Mux.scala 80:57]
  wire  _T_160_3 = _T_159 ? _T_618 : _T_158_3; // @[Mux.scala 80:57]
  wire  _T_162_3 = _T_161 ? _T_679 : _T_160_3; // @[Mux.scala 80:57]
  wire  _T_164_3 = _T_163 ? _T_740 : _T_162_3; // @[Mux.scala 80:57]
  wire  _T_166_3 = _T_165 ? _T_801 : _T_164_3; // @[Mux.scala 80:57]
  wire  _T_168_3 = _T_167 ? _T_862 : _T_166_3; // @[Mux.scala 80:57]
  wire  _T_170_3 = _T_169 ? _T_923 : _T_168_3; // @[Mux.scala 80:57]
  wire  _T_172_3 = _T_171 ? _T_984 : _T_170_3; // @[Mux.scala 80:57]
  wire  _T_174_3 = _T_173 ? _T_1045 : _T_172_3; // @[Mux.scala 80:57]
  wire  _T_176_3 = _T_175 ? _T_1106 : _T_174_3; // @[Mux.scala 80:57]
  wire  _T_178_3 = _T_177 ? _T_1167 : _T_176_3; // @[Mux.scala 80:57]
  wire  _T_180_3 = _T_179 ? _T_1228 : _T_178_3; // @[Mux.scala 80:57]
  wire  _T_182_3 = _T_181 ? _T_1289 : _T_180_3; // @[Mux.scala 80:57]
  wire  _T_184_3 = _T_183 ? _T_1350 : _T_182_3; // @[Mux.scala 80:57]
  wire  _T_186_3 = _T_185 ? _T_1411 : _T_184_3; // @[Mux.scala 80:57]
  wire  _T_188_3 = _T_187 ? _T_1472 : _T_186_3; // @[Mux.scala 80:57]
  wire  _T_190_3 = _T_189 ? _T_1533 : _T_188_3; // @[Mux.scala 80:57]
  wire  _T_192_3 = _T_191 ? _T_1594 : _T_190_3; // @[Mux.scala 80:57]
  wire  _T_194_3 = _T_193 ? _T_1655 : _T_192_3; // @[Mux.scala 80:57]
  wire  _T_196_3 = _T_195 ? _T_1716 : _T_194_3; // @[Mux.scala 80:57]
  wire  _T_198_3 = _T_197 ? _T_1777 : _T_196_3; // @[Mux.scala 80:57]
  wire  _T_200_3 = _T_199 ? _T_1838 : _T_198_3; // @[Mux.scala 80:57]
  wire  _T_202_3 = _T_201 ? _T_1899 : _T_200_3; // @[Mux.scala 80:57]
  wire  _T_204_3 = _T_203 ? _T_1960 : _T_202_3; // @[Mux.scala 80:57]
  wire  _T_206_3 = _T_205 ? _T_2021 : _T_204_3; // @[Mux.scala 80:57]
  wire  _T_208_3 = _T_207 ? _T_2082 : _T_206_3; // @[Mux.scala 80:57]
  wire  _T_210_3 = _T_209 ? _T_2143 : _T_208_3; // @[Mux.scala 80:57]
  wire  _T_212_3 = _T_211 ? _T_2204 : _T_210_3; // @[Mux.scala 80:57]
  wire  _T_214_3 = _T_213 ? _T_2265 : _T_212_3; // @[Mux.scala 80:57]
  wire  _T_216_3 = _T_215 ? _T_2326 : _T_214_3; // @[Mux.scala 80:57]
  wire  _T_218_3 = _T_217 ? _T_2387 : _T_216_3; // @[Mux.scala 80:57]
  wire  _T_220_3 = _T_219 ? _T_2448 : _T_218_3; // @[Mux.scala 80:57]
  wire  _T_222_3 = _T_221 ? _T_2509 : _T_220_3; // @[Mux.scala 80:57]
  wire  _T_224_3 = _T_223 ? _T_2570 : _T_222_3; // @[Mux.scala 80:57]
  wire  _T_226_3 = _T_225 ? _T_2631 : _T_224_3; // @[Mux.scala 80:57]
  wire  _T_228_3 = _T_227 ? _T_2692 : _T_226_3; // @[Mux.scala 80:57]
  wire  _T_230_3 = _T_229 ? _T_2753 : _T_228_3; // @[Mux.scala 80:57]
  wire  _T_232_3 = _T_231 ? _T_2814 : _T_230_3; // @[Mux.scala 80:57]
  wire  _T_234_3 = _T_233 ? _T_2875 : _T_232_3; // @[Mux.scala 80:57]
  wire  _T_236_3 = _T_235 ? _T_2936 : _T_234_3; // @[Mux.scala 80:57]
  wire  _T_238_3 = _T_237 ? _T_2997 : _T_236_3; // @[Mux.scala 80:57]
  wire  _T_240_3 = _T_239 ? _T_3058 : _T_238_3; // @[Mux.scala 80:57]
  wire  _T_242_3 = _T_241 ? _T_3119 : _T_240_3; // @[Mux.scala 80:57]
  wire  _T_244_3 = _T_243 ? _T_3180 : _T_242_3; // @[Mux.scala 80:57]
  wire  _T_246_3 = _T_245 ? _T_3241 : _T_244_3; // @[Mux.scala 80:57]
  wire  _T_248_3 = _T_247 ? _T_3302 : _T_246_3; // @[Mux.scala 80:57]
  wire  _T_250_3 = _T_249 ? _T_3363 : _T_248_3; // @[Mux.scala 80:57]
  wire  _T_252_3 = _T_251 ? _T_3424 : _T_250_3; // @[Mux.scala 80:57]
  wire  _T_254_3 = _T_253 ? _T_3485 : _T_252_3; // @[Mux.scala 80:57]
  wire  _T_256_3 = _T_255 ? _T_3546 : _T_254_3; // @[Mux.scala 80:57]
  wire  _T_258_3 = _T_257 ? _T_3607 : _T_256_3; // @[Mux.scala 80:57]
  wire  _T_260_3 = _T_259 ? _T_3668 : _T_258_3; // @[Mux.scala 80:57]
  wire  _T_262_3 = _T_261 ? _T_3729 : _T_260_3; // @[Mux.scala 80:57]
  wire  _T_264_3 = _T_263 ? _T_3790 : _T_262_3; // @[Mux.scala 80:57]
  wire  _T_266_3 = _T_265 ? _T_3851 : _T_264_3; // @[Mux.scala 80:57]
  wire  _T_268_3 = _T_267 ? _T_3912 : _T_266_3; // @[Mux.scala 80:57]
  wire  _T_270_3 = _T_269 ? _T_3973 : _T_268_3; // @[Mux.scala 80:57]
  wire  _T_272_3 = _T_271 ? _T_4034 : _T_270_3; // @[Mux.scala 80:57]
  wire  _T_274_3 = _T_273 ? _T_4095 : _T_272_3; // @[Mux.scala 80:57]
  wire  _T_276_3 = _T_275 ? _T_4156 : _T_274_3; // @[Mux.scala 80:57]
  wire  _T_278_3 = _T_277 ? _T_4217 : _T_276_3; // @[Mux.scala 80:57]
  wire  _T_280_3 = _T_279 ? _T_4278 : _T_278_3; // @[Mux.scala 80:57]
  wire  _T_282_3 = _T_281 ? _T_4339 : _T_280_3; // @[Mux.scala 80:57]
  reg [21:0] _T_4331; // @[Reg.scala 27:20]
  reg [21:0] _T_4270; // @[Reg.scala 27:20]
  reg [21:0] _T_4209; // @[Reg.scala 27:20]
  reg [21:0] _T_4148; // @[Reg.scala 27:20]
  reg [21:0] _T_4087; // @[Reg.scala 27:20]
  reg [21:0] _T_4026; // @[Reg.scala 27:20]
  reg [21:0] _T_3965; // @[Reg.scala 27:20]
  reg [21:0] _T_3904; // @[Reg.scala 27:20]
  reg [21:0] _T_3843; // @[Reg.scala 27:20]
  reg [21:0] _T_3782; // @[Reg.scala 27:20]
  reg [21:0] _T_3721; // @[Reg.scala 27:20]
  reg [21:0] _T_3660; // @[Reg.scala 27:20]
  reg [21:0] _T_3599; // @[Reg.scala 27:20]
  reg [21:0] _T_3538; // @[Reg.scala 27:20]
  reg [21:0] _T_3477; // @[Reg.scala 27:20]
  reg [21:0] _T_3416; // @[Reg.scala 27:20]
  reg [21:0] _T_3355; // @[Reg.scala 27:20]
  reg [21:0] _T_3294; // @[Reg.scala 27:20]
  reg [21:0] _T_3233; // @[Reg.scala 27:20]
  reg [21:0] _T_3172; // @[Reg.scala 27:20]
  reg [21:0] _T_3111; // @[Reg.scala 27:20]
  reg [21:0] _T_3050; // @[Reg.scala 27:20]
  reg [21:0] _T_2989; // @[Reg.scala 27:20]
  reg [21:0] _T_2928; // @[Reg.scala 27:20]
  reg [21:0] _T_2867; // @[Reg.scala 27:20]
  reg [21:0] _T_2806; // @[Reg.scala 27:20]
  reg [21:0] _T_2745; // @[Reg.scala 27:20]
  reg [21:0] _T_2684; // @[Reg.scala 27:20]
  reg [21:0] _T_2623; // @[Reg.scala 27:20]
  reg [21:0] _T_2562; // @[Reg.scala 27:20]
  reg [21:0] _T_2501; // @[Reg.scala 27:20]
  reg [21:0] _T_2440; // @[Reg.scala 27:20]
  reg [21:0] _T_2379; // @[Reg.scala 27:20]
  reg [21:0] _T_2318; // @[Reg.scala 27:20]
  reg [21:0] _T_2257; // @[Reg.scala 27:20]
  reg [21:0] _T_2196; // @[Reg.scala 27:20]
  reg [21:0] _T_2135; // @[Reg.scala 27:20]
  reg [21:0] _T_2074; // @[Reg.scala 27:20]
  reg [21:0] _T_2013; // @[Reg.scala 27:20]
  reg [21:0] _T_1952; // @[Reg.scala 27:20]
  reg [21:0] _T_1891; // @[Reg.scala 27:20]
  reg [21:0] _T_1830; // @[Reg.scala 27:20]
  reg [21:0] _T_1769; // @[Reg.scala 27:20]
  reg [21:0] _T_1708; // @[Reg.scala 27:20]
  reg [21:0] _T_1647; // @[Reg.scala 27:20]
  reg [21:0] _T_1586; // @[Reg.scala 27:20]
  reg [21:0] _T_1525; // @[Reg.scala 27:20]
  reg [21:0] _T_1464; // @[Reg.scala 27:20]
  reg [21:0] _T_1403; // @[Reg.scala 27:20]
  reg [21:0] _T_1342; // @[Reg.scala 27:20]
  reg [21:0] _T_1281; // @[Reg.scala 27:20]
  reg [21:0] _T_1220; // @[Reg.scala 27:20]
  reg [21:0] _T_1159; // @[Reg.scala 27:20]
  reg [21:0] _T_1098; // @[Reg.scala 27:20]
  reg [21:0] _T_1037; // @[Reg.scala 27:20]
  reg [21:0] _T_976; // @[Reg.scala 27:20]
  reg [21:0] _T_915; // @[Reg.scala 27:20]
  reg [21:0] _T_854; // @[Reg.scala 27:20]
  reg [21:0] _T_793; // @[Reg.scala 27:20]
  reg [21:0] _T_732; // @[Reg.scala 27:20]
  reg [21:0] _T_671; // @[Reg.scala 27:20]
  reg [21:0] _T_610; // @[Reg.scala 27:20]
  reg [21:0] _T_549; // @[Reg.scala 27:20]
  reg [21:0] _T_488; // @[Reg.scala 27:20]
  wire [21:0] _T_32_3 = _T_157 ? _T_549 : _T_488; // @[Mux.scala 80:57]
  wire [21:0] _T_34_3 = _T_159 ? _T_610 : _T_32_3; // @[Mux.scala 80:57]
  wire [21:0] _T_36_3 = _T_161 ? _T_671 : _T_34_3; // @[Mux.scala 80:57]
  wire [21:0] _T_38_3 = _T_163 ? _T_732 : _T_36_3; // @[Mux.scala 80:57]
  wire [21:0] _T_40_3 = _T_165 ? _T_793 : _T_38_3; // @[Mux.scala 80:57]
  wire [21:0] _T_42_3 = _T_167 ? _T_854 : _T_40_3; // @[Mux.scala 80:57]
  wire [21:0] _T_44_3 = _T_169 ? _T_915 : _T_42_3; // @[Mux.scala 80:57]
  wire [21:0] _T_46_3 = _T_171 ? _T_976 : _T_44_3; // @[Mux.scala 80:57]
  wire [21:0] _T_48_3 = _T_173 ? _T_1037 : _T_46_3; // @[Mux.scala 80:57]
  wire [21:0] _T_50_3 = _T_175 ? _T_1098 : _T_48_3; // @[Mux.scala 80:57]
  wire [21:0] _T_52_3 = _T_177 ? _T_1159 : _T_50_3; // @[Mux.scala 80:57]
  wire [21:0] _T_54_3 = _T_179 ? _T_1220 : _T_52_3; // @[Mux.scala 80:57]
  wire [21:0] _T_56_3 = _T_181 ? _T_1281 : _T_54_3; // @[Mux.scala 80:57]
  wire [21:0] _T_58_3 = _T_183 ? _T_1342 : _T_56_3; // @[Mux.scala 80:57]
  wire [21:0] _T_60_3 = _T_185 ? _T_1403 : _T_58_3; // @[Mux.scala 80:57]
  wire [21:0] _T_62_3 = _T_187 ? _T_1464 : _T_60_3; // @[Mux.scala 80:57]
  wire [21:0] _T_64_3 = _T_189 ? _T_1525 : _T_62_3; // @[Mux.scala 80:57]
  wire [21:0] _T_66_3 = _T_191 ? _T_1586 : _T_64_3; // @[Mux.scala 80:57]
  wire [21:0] _T_68_3 = _T_193 ? _T_1647 : _T_66_3; // @[Mux.scala 80:57]
  wire [21:0] _T_70_3 = _T_195 ? _T_1708 : _T_68_3; // @[Mux.scala 80:57]
  wire [21:0] _T_72_3 = _T_197 ? _T_1769 : _T_70_3; // @[Mux.scala 80:57]
  wire [21:0] _T_74_3 = _T_199 ? _T_1830 : _T_72_3; // @[Mux.scala 80:57]
  wire [21:0] _T_76_3 = _T_201 ? _T_1891 : _T_74_3; // @[Mux.scala 80:57]
  wire [21:0] _T_78_3 = _T_203 ? _T_1952 : _T_76_3; // @[Mux.scala 80:57]
  wire [21:0] _T_80_3 = _T_205 ? _T_2013 : _T_78_3; // @[Mux.scala 80:57]
  wire [21:0] _T_82_3 = _T_207 ? _T_2074 : _T_80_3; // @[Mux.scala 80:57]
  wire [21:0] _T_84_3 = _T_209 ? _T_2135 : _T_82_3; // @[Mux.scala 80:57]
  wire [21:0] _T_86_3 = _T_211 ? _T_2196 : _T_84_3; // @[Mux.scala 80:57]
  wire [21:0] _T_88_3 = _T_213 ? _T_2257 : _T_86_3; // @[Mux.scala 80:57]
  wire [21:0] _T_90_3 = _T_215 ? _T_2318 : _T_88_3; // @[Mux.scala 80:57]
  wire [21:0] _T_92_3 = _T_217 ? _T_2379 : _T_90_3; // @[Mux.scala 80:57]
  wire [21:0] _T_94_3 = _T_219 ? _T_2440 : _T_92_3; // @[Mux.scala 80:57]
  wire [21:0] _T_96_3 = _T_221 ? _T_2501 : _T_94_3; // @[Mux.scala 80:57]
  wire [21:0] _T_98_3 = _T_223 ? _T_2562 : _T_96_3; // @[Mux.scala 80:57]
  wire [21:0] _T_100_3 = _T_225 ? _T_2623 : _T_98_3; // @[Mux.scala 80:57]
  wire [21:0] _T_102_3 = _T_227 ? _T_2684 : _T_100_3; // @[Mux.scala 80:57]
  wire [21:0] _T_104_3 = _T_229 ? _T_2745 : _T_102_3; // @[Mux.scala 80:57]
  wire [21:0] _T_106_3 = _T_231 ? _T_2806 : _T_104_3; // @[Mux.scala 80:57]
  wire [21:0] _T_108_3 = _T_233 ? _T_2867 : _T_106_3; // @[Mux.scala 80:57]
  wire [21:0] _T_110_3 = _T_235 ? _T_2928 : _T_108_3; // @[Mux.scala 80:57]
  wire [21:0] _T_112_3 = _T_237 ? _T_2989 : _T_110_3; // @[Mux.scala 80:57]
  wire [21:0] _T_114_3 = _T_239 ? _T_3050 : _T_112_3; // @[Mux.scala 80:57]
  wire [21:0] _T_116_3 = _T_241 ? _T_3111 : _T_114_3; // @[Mux.scala 80:57]
  wire [21:0] _T_118_3 = _T_243 ? _T_3172 : _T_116_3; // @[Mux.scala 80:57]
  wire [21:0] _T_120_3 = _T_245 ? _T_3233 : _T_118_3; // @[Mux.scala 80:57]
  wire [21:0] _T_122_3 = _T_247 ? _T_3294 : _T_120_3; // @[Mux.scala 80:57]
  wire [21:0] _T_124_3 = _T_249 ? _T_3355 : _T_122_3; // @[Mux.scala 80:57]
  wire [21:0] _T_126_3 = _T_251 ? _T_3416 : _T_124_3; // @[Mux.scala 80:57]
  wire [21:0] _T_128_3 = _T_253 ? _T_3477 : _T_126_3; // @[Mux.scala 80:57]
  wire [21:0] _T_130_3 = _T_255 ? _T_3538 : _T_128_3; // @[Mux.scala 80:57]
  wire [21:0] _T_132_3 = _T_257 ? _T_3599 : _T_130_3; // @[Mux.scala 80:57]
  wire [21:0] _T_134_3 = _T_259 ? _T_3660 : _T_132_3; // @[Mux.scala 80:57]
  wire [21:0] _T_136_3 = _T_261 ? _T_3721 : _T_134_3; // @[Mux.scala 80:57]
  wire [21:0] _T_138_3 = _T_263 ? _T_3782 : _T_136_3; // @[Mux.scala 80:57]
  wire [21:0] _T_140_3 = _T_265 ? _T_3843 : _T_138_3; // @[Mux.scala 80:57]
  wire [21:0] _T_142_3 = _T_267 ? _T_3904 : _T_140_3; // @[Mux.scala 80:57]
  wire [21:0] _T_144_3 = _T_269 ? _T_3965 : _T_142_3; // @[Mux.scala 80:57]
  wire [21:0] _T_146_3 = _T_271 ? _T_4026 : _T_144_3; // @[Mux.scala 80:57]
  wire [21:0] _T_148_3 = _T_273 ? _T_4087 : _T_146_3; // @[Mux.scala 80:57]
  wire [21:0] _T_150_3 = _T_275 ? _T_4148 : _T_148_3; // @[Mux.scala 80:57]
  wire [21:0] _T_152_3 = _T_277 ? _T_4209 : _T_150_3; // @[Mux.scala 80:57]
  wire [21:0] _T_154_3 = _T_279 ? _T_4270 : _T_152_3; // @[Mux.scala 80:57]
  wire [21:0] _T_156_3 = _T_281 ? _T_4331 : _T_154_3; // @[Mux.scala 80:57]
  wire  _T_289 = _T_156_3 == io_cacheIn_addr[31:10]; // @[Cache.scala 772:78]
  wire  _T_290 = _T_282_3 & _T_289; // @[Cache.scala 772:62]
  wire  _T_294 = _T_293 | _T_290; // @[Cache.scala 773:51]
  wire  _T_14 = 3'h0 == _T_4; // @[Mux.scala 80:60]
  wire  _T_16 = 3'h1 == _T_4; // @[Mux.scala 80:60]
  wire  _T_18 = 3'h2 == _T_4; // @[Mux.scala 80:60]
  wire  _T_20 = 3'h3 == _T_4; // @[Mux.scala 80:60]
  wire  _T_22 = 3'h4 == _T_4; // @[Mux.scala 80:60]
  wire  _T_24 = _T_4 == 3'h0; // @[Cache.scala 742:29]
  wire  _T_25 = _T_4 == 3'h1; // @[Cache.scala 743:29]
  wire  _T_26 = _T_4 == 3'h2; // @[Cache.scala 744:29]
  wire  _T_27 = _T_4 == 3'h3; // @[Cache.scala 745:30]
  wire  _T_28 = _T_4 == 3'h4; // @[Cache.scala 746:30]
  wire [127:0] _T_295 = _T_284 ? io_SRAMIO_0_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _T_296 = _T_286 ? io_SRAMIO_1_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _T_297 = _T_288 ? io_SRAMIO_2_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _T_298 = _T_290 ? io_SRAMIO_3_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _T_299 = _T_295 | _T_296; // @[Mux.scala 27:72]
  wire [127:0] _T_300 = _T_299 | _T_297; // @[Mux.scala 27:72]
  wire [127:0] _T_301 = _T_300 | _T_298; // @[Mux.scala 27:72]
  reg [1:0] _T_501; // @[Reg.scala 27:20]
  reg [1:0] _T_440; // @[Reg.scala 27:20]
  wire [1:0] _T_309 = _T_157 ? _T_501 : _T_440; // @[Mux.scala 80:57]
  reg [1:0] _T_562; // @[Reg.scala 27:20]
  wire [1:0] _T_311 = _T_159 ? _T_562 : _T_309; // @[Mux.scala 80:57]
  reg [1:0] _T_623; // @[Reg.scala 27:20]
  wire [1:0] _T_313 = _T_161 ? _T_623 : _T_311; // @[Mux.scala 80:57]
  reg [1:0] _T_684; // @[Reg.scala 27:20]
  wire [1:0] _T_315 = _T_163 ? _T_684 : _T_313; // @[Mux.scala 80:57]
  reg [1:0] _T_745; // @[Reg.scala 27:20]
  wire [1:0] _T_317 = _T_165 ? _T_745 : _T_315; // @[Mux.scala 80:57]
  reg [1:0] _T_806; // @[Reg.scala 27:20]
  wire [1:0] _T_319 = _T_167 ? _T_806 : _T_317; // @[Mux.scala 80:57]
  reg [1:0] _T_867; // @[Reg.scala 27:20]
  wire [1:0] _T_321 = _T_169 ? _T_867 : _T_319; // @[Mux.scala 80:57]
  reg [1:0] _T_928; // @[Reg.scala 27:20]
  wire [1:0] _T_323 = _T_171 ? _T_928 : _T_321; // @[Mux.scala 80:57]
  reg [1:0] _T_989; // @[Reg.scala 27:20]
  wire [1:0] _T_325 = _T_173 ? _T_989 : _T_323; // @[Mux.scala 80:57]
  reg [1:0] _T_1050; // @[Reg.scala 27:20]
  wire [1:0] _T_327 = _T_175 ? _T_1050 : _T_325; // @[Mux.scala 80:57]
  reg [1:0] _T_1111; // @[Reg.scala 27:20]
  wire [1:0] _T_329 = _T_177 ? _T_1111 : _T_327; // @[Mux.scala 80:57]
  reg [1:0] _T_1172; // @[Reg.scala 27:20]
  wire [1:0] _T_331 = _T_179 ? _T_1172 : _T_329; // @[Mux.scala 80:57]
  reg [1:0] _T_1233; // @[Reg.scala 27:20]
  wire [1:0] _T_333 = _T_181 ? _T_1233 : _T_331; // @[Mux.scala 80:57]
  reg [1:0] _T_1294; // @[Reg.scala 27:20]
  wire [1:0] _T_335 = _T_183 ? _T_1294 : _T_333; // @[Mux.scala 80:57]
  reg [1:0] _T_1355; // @[Reg.scala 27:20]
  wire [1:0] _T_337 = _T_185 ? _T_1355 : _T_335; // @[Mux.scala 80:57]
  reg [1:0] _T_1416; // @[Reg.scala 27:20]
  wire [1:0] _T_339 = _T_187 ? _T_1416 : _T_337; // @[Mux.scala 80:57]
  reg [1:0] _T_1477; // @[Reg.scala 27:20]
  wire [1:0] _T_341 = _T_189 ? _T_1477 : _T_339; // @[Mux.scala 80:57]
  reg [1:0] _T_1538; // @[Reg.scala 27:20]
  wire [1:0] _T_343 = _T_191 ? _T_1538 : _T_341; // @[Mux.scala 80:57]
  reg [1:0] _T_1599; // @[Reg.scala 27:20]
  wire [1:0] _T_345 = _T_193 ? _T_1599 : _T_343; // @[Mux.scala 80:57]
  reg [1:0] _T_1660; // @[Reg.scala 27:20]
  wire [1:0] _T_347 = _T_195 ? _T_1660 : _T_345; // @[Mux.scala 80:57]
  reg [1:0] _T_1721; // @[Reg.scala 27:20]
  wire [1:0] _T_349 = _T_197 ? _T_1721 : _T_347; // @[Mux.scala 80:57]
  reg [1:0] _T_1782; // @[Reg.scala 27:20]
  wire [1:0] _T_351 = _T_199 ? _T_1782 : _T_349; // @[Mux.scala 80:57]
  reg [1:0] _T_1843; // @[Reg.scala 27:20]
  wire [1:0] _T_353 = _T_201 ? _T_1843 : _T_351; // @[Mux.scala 80:57]
  reg [1:0] _T_1904; // @[Reg.scala 27:20]
  wire [1:0] _T_355 = _T_203 ? _T_1904 : _T_353; // @[Mux.scala 80:57]
  reg [1:0] _T_1965; // @[Reg.scala 27:20]
  wire [1:0] _T_357 = _T_205 ? _T_1965 : _T_355; // @[Mux.scala 80:57]
  reg [1:0] _T_2026; // @[Reg.scala 27:20]
  wire [1:0] _T_359 = _T_207 ? _T_2026 : _T_357; // @[Mux.scala 80:57]
  reg [1:0] _T_2087; // @[Reg.scala 27:20]
  wire [1:0] _T_361 = _T_209 ? _T_2087 : _T_359; // @[Mux.scala 80:57]
  reg [1:0] _T_2148; // @[Reg.scala 27:20]
  wire [1:0] _T_363 = _T_211 ? _T_2148 : _T_361; // @[Mux.scala 80:57]
  reg [1:0] _T_2209; // @[Reg.scala 27:20]
  wire [1:0] _T_365 = _T_213 ? _T_2209 : _T_363; // @[Mux.scala 80:57]
  reg [1:0] _T_2270; // @[Reg.scala 27:20]
  wire [1:0] _T_367 = _T_215 ? _T_2270 : _T_365; // @[Mux.scala 80:57]
  reg [1:0] _T_2331; // @[Reg.scala 27:20]
  wire [1:0] _T_369 = _T_217 ? _T_2331 : _T_367; // @[Mux.scala 80:57]
  reg [1:0] _T_2392; // @[Reg.scala 27:20]
  wire [1:0] _T_371 = _T_219 ? _T_2392 : _T_369; // @[Mux.scala 80:57]
  reg [1:0] _T_2453; // @[Reg.scala 27:20]
  wire [1:0] _T_373 = _T_221 ? _T_2453 : _T_371; // @[Mux.scala 80:57]
  reg [1:0] _T_2514; // @[Reg.scala 27:20]
  wire [1:0] _T_375 = _T_223 ? _T_2514 : _T_373; // @[Mux.scala 80:57]
  reg [1:0] _T_2575; // @[Reg.scala 27:20]
  wire [1:0] _T_377 = _T_225 ? _T_2575 : _T_375; // @[Mux.scala 80:57]
  reg [1:0] _T_2636; // @[Reg.scala 27:20]
  wire [1:0] _T_379 = _T_227 ? _T_2636 : _T_377; // @[Mux.scala 80:57]
  reg [1:0] _T_2697; // @[Reg.scala 27:20]
  wire [1:0] _T_381 = _T_229 ? _T_2697 : _T_379; // @[Mux.scala 80:57]
  reg [1:0] _T_2758; // @[Reg.scala 27:20]
  wire [1:0] _T_383 = _T_231 ? _T_2758 : _T_381; // @[Mux.scala 80:57]
  reg [1:0] _T_2819; // @[Reg.scala 27:20]
  wire [1:0] _T_385 = _T_233 ? _T_2819 : _T_383; // @[Mux.scala 80:57]
  reg [1:0] _T_2880; // @[Reg.scala 27:20]
  wire [1:0] _T_387 = _T_235 ? _T_2880 : _T_385; // @[Mux.scala 80:57]
  reg [1:0] _T_2941; // @[Reg.scala 27:20]
  wire [1:0] _T_389 = _T_237 ? _T_2941 : _T_387; // @[Mux.scala 80:57]
  reg [1:0] _T_3002; // @[Reg.scala 27:20]
  wire [1:0] _T_391 = _T_239 ? _T_3002 : _T_389; // @[Mux.scala 80:57]
  reg [1:0] _T_3063; // @[Reg.scala 27:20]
  wire [1:0] _T_393 = _T_241 ? _T_3063 : _T_391; // @[Mux.scala 80:57]
  reg [1:0] _T_3124; // @[Reg.scala 27:20]
  wire [1:0] _T_395 = _T_243 ? _T_3124 : _T_393; // @[Mux.scala 80:57]
  reg [1:0] _T_3185; // @[Reg.scala 27:20]
  wire [1:0] _T_397 = _T_245 ? _T_3185 : _T_395; // @[Mux.scala 80:57]
  reg [1:0] _T_3246; // @[Reg.scala 27:20]
  wire [1:0] _T_399 = _T_247 ? _T_3246 : _T_397; // @[Mux.scala 80:57]
  reg [1:0] _T_3307; // @[Reg.scala 27:20]
  wire [1:0] _T_401 = _T_249 ? _T_3307 : _T_399; // @[Mux.scala 80:57]
  reg [1:0] _T_3368; // @[Reg.scala 27:20]
  wire [1:0] _T_403 = _T_251 ? _T_3368 : _T_401; // @[Mux.scala 80:57]
  reg [1:0] _T_3429; // @[Reg.scala 27:20]
  wire [1:0] _T_405 = _T_253 ? _T_3429 : _T_403; // @[Mux.scala 80:57]
  reg [1:0] _T_3490; // @[Reg.scala 27:20]
  wire [1:0] _T_407 = _T_255 ? _T_3490 : _T_405; // @[Mux.scala 80:57]
  reg [1:0] _T_3551; // @[Reg.scala 27:20]
  wire [1:0] _T_409 = _T_257 ? _T_3551 : _T_407; // @[Mux.scala 80:57]
  reg [1:0] _T_3612; // @[Reg.scala 27:20]
  wire [1:0] _T_411 = _T_259 ? _T_3612 : _T_409; // @[Mux.scala 80:57]
  reg [1:0] _T_3673; // @[Reg.scala 27:20]
  wire [1:0] _T_413 = _T_261 ? _T_3673 : _T_411; // @[Mux.scala 80:57]
  reg [1:0] _T_3734; // @[Reg.scala 27:20]
  wire [1:0] _T_415 = _T_263 ? _T_3734 : _T_413; // @[Mux.scala 80:57]
  reg [1:0] _T_3795; // @[Reg.scala 27:20]
  wire [1:0] _T_417 = _T_265 ? _T_3795 : _T_415; // @[Mux.scala 80:57]
  reg [1:0] _T_3856; // @[Reg.scala 27:20]
  wire [1:0] _T_419 = _T_267 ? _T_3856 : _T_417; // @[Mux.scala 80:57]
  reg [1:0] _T_3917; // @[Reg.scala 27:20]
  wire [1:0] _T_421 = _T_269 ? _T_3917 : _T_419; // @[Mux.scala 80:57]
  reg [1:0] _T_3978; // @[Reg.scala 27:20]
  wire [1:0] _T_423 = _T_271 ? _T_3978 : _T_421; // @[Mux.scala 80:57]
  reg [1:0] _T_4039; // @[Reg.scala 27:20]
  wire [1:0] _T_425 = _T_273 ? _T_4039 : _T_423; // @[Mux.scala 80:57]
  reg [1:0] _T_4100; // @[Reg.scala 27:20]
  wire [1:0] _T_427 = _T_275 ? _T_4100 : _T_425; // @[Mux.scala 80:57]
  reg [1:0] _T_4161; // @[Reg.scala 27:20]
  wire [1:0] _T_429 = _T_277 ? _T_4161 : _T_427; // @[Mux.scala 80:57]
  reg [1:0] _T_4222; // @[Reg.scala 27:20]
  wire [1:0] _T_431 = _T_279 ? _T_4222 : _T_429; // @[Mux.scala 80:57]
  reg [1:0] _T_4283; // @[Reg.scala 27:20]
  wire [1:0] _T_433 = _T_281 ? _T_4283 : _T_431; // @[Mux.scala 80:57]
  wire [1:0] _T_437 = _T_440 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_438 = 6'h0 == io_cacheIn_addr[9:4]; // @[Cache.scala 824:37]
  wire  _T_439 = io_cacheOut_r_last_i & _T_438; // @[Cache.scala 824:30]
  wire  _T_443 = _T_440 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_444 = _T_439 & _T_443; // @[Cache.scala 827:89]
  wire  _T_445 = _T_444 & _T_25; // @[Cache.scala 827:116]
  wire  _T_448 = reset | updataICache; // @[Cache.scala 828:34]
  wire  _GEN_2 = _T_445 | _T_454; // @[Reg.scala 28:19]
  wire  _T_457 = _T_440 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_458 = _T_439 & _T_457; // @[Cache.scala 827:89]
  wire  _T_459 = _T_458 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_4 = _T_459 | _T_468; // @[Reg.scala 28:19]
  wire  _T_471 = _T_440 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_472 = _T_439 & _T_471; // @[Cache.scala 827:89]
  wire  _T_473 = _T_472 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_6 = _T_473 | _T_482; // @[Reg.scala 28:19]
  wire  _T_485 = _T_440 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_486 = _T_439 & _T_485; // @[Cache.scala 827:89]
  wire  _T_487 = _T_486 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_8 = _T_487 | _T_496; // @[Reg.scala 28:19]
  wire [1:0] _T_498 = _T_501 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_500 = io_cacheOut_r_last_i & _T_157; // @[Cache.scala 824:30]
  wire  _T_504 = _T_501 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_505 = _T_500 & _T_504; // @[Cache.scala 827:89]
  wire  _T_506 = _T_505 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_11 = _T_506 | _T_515; // @[Reg.scala 28:19]
  wire  _T_518 = _T_501 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_519 = _T_500 & _T_518; // @[Cache.scala 827:89]
  wire  _T_520 = _T_519 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_13 = _T_520 | _T_529; // @[Reg.scala 28:19]
  wire  _T_532 = _T_501 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_533 = _T_500 & _T_532; // @[Cache.scala 827:89]
  wire  _T_534 = _T_533 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_15 = _T_534 | _T_543; // @[Reg.scala 28:19]
  wire  _T_546 = _T_501 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_547 = _T_500 & _T_546; // @[Cache.scala 827:89]
  wire  _T_548 = _T_547 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_17 = _T_548 | _T_557; // @[Reg.scala 28:19]
  wire [1:0] _T_559 = _T_562 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_561 = io_cacheOut_r_last_i & _T_159; // @[Cache.scala 824:30]
  wire  _T_565 = _T_562 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_566 = _T_561 & _T_565; // @[Cache.scala 827:89]
  wire  _T_567 = _T_566 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_20 = _T_567 | _T_576; // @[Reg.scala 28:19]
  wire  _T_579 = _T_562 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_580 = _T_561 & _T_579; // @[Cache.scala 827:89]
  wire  _T_581 = _T_580 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_22 = _T_581 | _T_590; // @[Reg.scala 28:19]
  wire  _T_593 = _T_562 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_594 = _T_561 & _T_593; // @[Cache.scala 827:89]
  wire  _T_595 = _T_594 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_24 = _T_595 | _T_604; // @[Reg.scala 28:19]
  wire  _T_607 = _T_562 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_608 = _T_561 & _T_607; // @[Cache.scala 827:89]
  wire  _T_609 = _T_608 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_26 = _T_609 | _T_618; // @[Reg.scala 28:19]
  wire [1:0] _T_620 = _T_623 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_622 = io_cacheOut_r_last_i & _T_161; // @[Cache.scala 824:30]
  wire  _T_626 = _T_623 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_627 = _T_622 & _T_626; // @[Cache.scala 827:89]
  wire  _T_628 = _T_627 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_29 = _T_628 | _T_637; // @[Reg.scala 28:19]
  wire  _T_640 = _T_623 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_641 = _T_622 & _T_640; // @[Cache.scala 827:89]
  wire  _T_642 = _T_641 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_31 = _T_642 | _T_651; // @[Reg.scala 28:19]
  wire  _T_654 = _T_623 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_655 = _T_622 & _T_654; // @[Cache.scala 827:89]
  wire  _T_656 = _T_655 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_33 = _T_656 | _T_665; // @[Reg.scala 28:19]
  wire  _T_668 = _T_623 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_669 = _T_622 & _T_668; // @[Cache.scala 827:89]
  wire  _T_670 = _T_669 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_35 = _T_670 | _T_679; // @[Reg.scala 28:19]
  wire [1:0] _T_681 = _T_684 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_683 = io_cacheOut_r_last_i & _T_163; // @[Cache.scala 824:30]
  wire  _T_687 = _T_684 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_688 = _T_683 & _T_687; // @[Cache.scala 827:89]
  wire  _T_689 = _T_688 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_38 = _T_689 | _T_698; // @[Reg.scala 28:19]
  wire  _T_701 = _T_684 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_702 = _T_683 & _T_701; // @[Cache.scala 827:89]
  wire  _T_703 = _T_702 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_40 = _T_703 | _T_712; // @[Reg.scala 28:19]
  wire  _T_715 = _T_684 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_716 = _T_683 & _T_715; // @[Cache.scala 827:89]
  wire  _T_717 = _T_716 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_42 = _T_717 | _T_726; // @[Reg.scala 28:19]
  wire  _T_729 = _T_684 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_730 = _T_683 & _T_729; // @[Cache.scala 827:89]
  wire  _T_731 = _T_730 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_44 = _T_731 | _T_740; // @[Reg.scala 28:19]
  wire [1:0] _T_742 = _T_745 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_744 = io_cacheOut_r_last_i & _T_165; // @[Cache.scala 824:30]
  wire  _T_748 = _T_745 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_749 = _T_744 & _T_748; // @[Cache.scala 827:89]
  wire  _T_750 = _T_749 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_47 = _T_750 | _T_759; // @[Reg.scala 28:19]
  wire  _T_762 = _T_745 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_763 = _T_744 & _T_762; // @[Cache.scala 827:89]
  wire  _T_764 = _T_763 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_49 = _T_764 | _T_773; // @[Reg.scala 28:19]
  wire  _T_776 = _T_745 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_777 = _T_744 & _T_776; // @[Cache.scala 827:89]
  wire  _T_778 = _T_777 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_51 = _T_778 | _T_787; // @[Reg.scala 28:19]
  wire  _T_790 = _T_745 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_791 = _T_744 & _T_790; // @[Cache.scala 827:89]
  wire  _T_792 = _T_791 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_53 = _T_792 | _T_801; // @[Reg.scala 28:19]
  wire [1:0] _T_803 = _T_806 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_805 = io_cacheOut_r_last_i & _T_167; // @[Cache.scala 824:30]
  wire  _T_809 = _T_806 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_810 = _T_805 & _T_809; // @[Cache.scala 827:89]
  wire  _T_811 = _T_810 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_56 = _T_811 | _T_820; // @[Reg.scala 28:19]
  wire  _T_823 = _T_806 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_824 = _T_805 & _T_823; // @[Cache.scala 827:89]
  wire  _T_825 = _T_824 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_58 = _T_825 | _T_834; // @[Reg.scala 28:19]
  wire  _T_837 = _T_806 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_838 = _T_805 & _T_837; // @[Cache.scala 827:89]
  wire  _T_839 = _T_838 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_60 = _T_839 | _T_848; // @[Reg.scala 28:19]
  wire  _T_851 = _T_806 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_852 = _T_805 & _T_851; // @[Cache.scala 827:89]
  wire  _T_853 = _T_852 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_62 = _T_853 | _T_862; // @[Reg.scala 28:19]
  wire [1:0] _T_864 = _T_867 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_866 = io_cacheOut_r_last_i & _T_169; // @[Cache.scala 824:30]
  wire  _T_870 = _T_867 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_871 = _T_866 & _T_870; // @[Cache.scala 827:89]
  wire  _T_872 = _T_871 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_65 = _T_872 | _T_881; // @[Reg.scala 28:19]
  wire  _T_884 = _T_867 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_885 = _T_866 & _T_884; // @[Cache.scala 827:89]
  wire  _T_886 = _T_885 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_67 = _T_886 | _T_895; // @[Reg.scala 28:19]
  wire  _T_898 = _T_867 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_899 = _T_866 & _T_898; // @[Cache.scala 827:89]
  wire  _T_900 = _T_899 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_69 = _T_900 | _T_909; // @[Reg.scala 28:19]
  wire  _T_912 = _T_867 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_913 = _T_866 & _T_912; // @[Cache.scala 827:89]
  wire  _T_914 = _T_913 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_71 = _T_914 | _T_923; // @[Reg.scala 28:19]
  wire [1:0] _T_925 = _T_928 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_927 = io_cacheOut_r_last_i & _T_171; // @[Cache.scala 824:30]
  wire  _T_931 = _T_928 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_932 = _T_927 & _T_931; // @[Cache.scala 827:89]
  wire  _T_933 = _T_932 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_74 = _T_933 | _T_942; // @[Reg.scala 28:19]
  wire  _T_945 = _T_928 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_946 = _T_927 & _T_945; // @[Cache.scala 827:89]
  wire  _T_947 = _T_946 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_76 = _T_947 | _T_956; // @[Reg.scala 28:19]
  wire  _T_959 = _T_928 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_960 = _T_927 & _T_959; // @[Cache.scala 827:89]
  wire  _T_961 = _T_960 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_78 = _T_961 | _T_970; // @[Reg.scala 28:19]
  wire  _T_973 = _T_928 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_974 = _T_927 & _T_973; // @[Cache.scala 827:89]
  wire  _T_975 = _T_974 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_80 = _T_975 | _T_984; // @[Reg.scala 28:19]
  wire [1:0] _T_986 = _T_989 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_988 = io_cacheOut_r_last_i & _T_173; // @[Cache.scala 824:30]
  wire  _T_992 = _T_989 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_993 = _T_988 & _T_992; // @[Cache.scala 827:89]
  wire  _T_994 = _T_993 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_83 = _T_994 | _T_1003; // @[Reg.scala 28:19]
  wire  _T_1006 = _T_989 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_1007 = _T_988 & _T_1006; // @[Cache.scala 827:89]
  wire  _T_1008 = _T_1007 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_85 = _T_1008 | _T_1017; // @[Reg.scala 28:19]
  wire  _T_1020 = _T_989 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_1021 = _T_988 & _T_1020; // @[Cache.scala 827:89]
  wire  _T_1022 = _T_1021 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_87 = _T_1022 | _T_1031; // @[Reg.scala 28:19]
  wire  _T_1034 = _T_989 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_1035 = _T_988 & _T_1034; // @[Cache.scala 827:89]
  wire  _T_1036 = _T_1035 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_89 = _T_1036 | _T_1045; // @[Reg.scala 28:19]
  wire [1:0] _T_1047 = _T_1050 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_1049 = io_cacheOut_r_last_i & _T_175; // @[Cache.scala 824:30]
  wire  _T_1053 = _T_1050 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_1054 = _T_1049 & _T_1053; // @[Cache.scala 827:89]
  wire  _T_1055 = _T_1054 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_92 = _T_1055 | _T_1064; // @[Reg.scala 28:19]
  wire  _T_1067 = _T_1050 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_1068 = _T_1049 & _T_1067; // @[Cache.scala 827:89]
  wire  _T_1069 = _T_1068 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_94 = _T_1069 | _T_1078; // @[Reg.scala 28:19]
  wire  _T_1081 = _T_1050 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_1082 = _T_1049 & _T_1081; // @[Cache.scala 827:89]
  wire  _T_1083 = _T_1082 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_96 = _T_1083 | _T_1092; // @[Reg.scala 28:19]
  wire  _T_1095 = _T_1050 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_1096 = _T_1049 & _T_1095; // @[Cache.scala 827:89]
  wire  _T_1097 = _T_1096 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_98 = _T_1097 | _T_1106; // @[Reg.scala 28:19]
  wire [1:0] _T_1108 = _T_1111 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_1110 = io_cacheOut_r_last_i & _T_177; // @[Cache.scala 824:30]
  wire  _T_1114 = _T_1111 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_1115 = _T_1110 & _T_1114; // @[Cache.scala 827:89]
  wire  _T_1116 = _T_1115 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_101 = _T_1116 | _T_1125; // @[Reg.scala 28:19]
  wire  _T_1128 = _T_1111 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_1129 = _T_1110 & _T_1128; // @[Cache.scala 827:89]
  wire  _T_1130 = _T_1129 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_103 = _T_1130 | _T_1139; // @[Reg.scala 28:19]
  wire  _T_1142 = _T_1111 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_1143 = _T_1110 & _T_1142; // @[Cache.scala 827:89]
  wire  _T_1144 = _T_1143 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_105 = _T_1144 | _T_1153; // @[Reg.scala 28:19]
  wire  _T_1156 = _T_1111 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_1157 = _T_1110 & _T_1156; // @[Cache.scala 827:89]
  wire  _T_1158 = _T_1157 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_107 = _T_1158 | _T_1167; // @[Reg.scala 28:19]
  wire [1:0] _T_1169 = _T_1172 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_1171 = io_cacheOut_r_last_i & _T_179; // @[Cache.scala 824:30]
  wire  _T_1175 = _T_1172 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_1176 = _T_1171 & _T_1175; // @[Cache.scala 827:89]
  wire  _T_1177 = _T_1176 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_110 = _T_1177 | _T_1186; // @[Reg.scala 28:19]
  wire  _T_1189 = _T_1172 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_1190 = _T_1171 & _T_1189; // @[Cache.scala 827:89]
  wire  _T_1191 = _T_1190 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_112 = _T_1191 | _T_1200; // @[Reg.scala 28:19]
  wire  _T_1203 = _T_1172 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_1204 = _T_1171 & _T_1203; // @[Cache.scala 827:89]
  wire  _T_1205 = _T_1204 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_114 = _T_1205 | _T_1214; // @[Reg.scala 28:19]
  wire  _T_1217 = _T_1172 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_1218 = _T_1171 & _T_1217; // @[Cache.scala 827:89]
  wire  _T_1219 = _T_1218 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_116 = _T_1219 | _T_1228; // @[Reg.scala 28:19]
  wire [1:0] _T_1230 = _T_1233 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_1232 = io_cacheOut_r_last_i & _T_181; // @[Cache.scala 824:30]
  wire  _T_1236 = _T_1233 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_1237 = _T_1232 & _T_1236; // @[Cache.scala 827:89]
  wire  _T_1238 = _T_1237 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_119 = _T_1238 | _T_1247; // @[Reg.scala 28:19]
  wire  _T_1250 = _T_1233 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_1251 = _T_1232 & _T_1250; // @[Cache.scala 827:89]
  wire  _T_1252 = _T_1251 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_121 = _T_1252 | _T_1261; // @[Reg.scala 28:19]
  wire  _T_1264 = _T_1233 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_1265 = _T_1232 & _T_1264; // @[Cache.scala 827:89]
  wire  _T_1266 = _T_1265 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_123 = _T_1266 | _T_1275; // @[Reg.scala 28:19]
  wire  _T_1278 = _T_1233 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_1279 = _T_1232 & _T_1278; // @[Cache.scala 827:89]
  wire  _T_1280 = _T_1279 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_125 = _T_1280 | _T_1289; // @[Reg.scala 28:19]
  wire [1:0] _T_1291 = _T_1294 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_1293 = io_cacheOut_r_last_i & _T_183; // @[Cache.scala 824:30]
  wire  _T_1297 = _T_1294 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_1298 = _T_1293 & _T_1297; // @[Cache.scala 827:89]
  wire  _T_1299 = _T_1298 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_128 = _T_1299 | _T_1308; // @[Reg.scala 28:19]
  wire  _T_1311 = _T_1294 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_1312 = _T_1293 & _T_1311; // @[Cache.scala 827:89]
  wire  _T_1313 = _T_1312 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_130 = _T_1313 | _T_1322; // @[Reg.scala 28:19]
  wire  _T_1325 = _T_1294 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_1326 = _T_1293 & _T_1325; // @[Cache.scala 827:89]
  wire  _T_1327 = _T_1326 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_132 = _T_1327 | _T_1336; // @[Reg.scala 28:19]
  wire  _T_1339 = _T_1294 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_1340 = _T_1293 & _T_1339; // @[Cache.scala 827:89]
  wire  _T_1341 = _T_1340 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_134 = _T_1341 | _T_1350; // @[Reg.scala 28:19]
  wire [1:0] _T_1352 = _T_1355 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_1354 = io_cacheOut_r_last_i & _T_185; // @[Cache.scala 824:30]
  wire  _T_1358 = _T_1355 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_1359 = _T_1354 & _T_1358; // @[Cache.scala 827:89]
  wire  _T_1360 = _T_1359 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_137 = _T_1360 | _T_1369; // @[Reg.scala 28:19]
  wire  _T_1372 = _T_1355 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_1373 = _T_1354 & _T_1372; // @[Cache.scala 827:89]
  wire  _T_1374 = _T_1373 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_139 = _T_1374 | _T_1383; // @[Reg.scala 28:19]
  wire  _T_1386 = _T_1355 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_1387 = _T_1354 & _T_1386; // @[Cache.scala 827:89]
  wire  _T_1388 = _T_1387 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_141 = _T_1388 | _T_1397; // @[Reg.scala 28:19]
  wire  _T_1400 = _T_1355 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_1401 = _T_1354 & _T_1400; // @[Cache.scala 827:89]
  wire  _T_1402 = _T_1401 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_143 = _T_1402 | _T_1411; // @[Reg.scala 28:19]
  wire [1:0] _T_1413 = _T_1416 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_1415 = io_cacheOut_r_last_i & _T_187; // @[Cache.scala 824:30]
  wire  _T_1419 = _T_1416 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_1420 = _T_1415 & _T_1419; // @[Cache.scala 827:89]
  wire  _T_1421 = _T_1420 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_146 = _T_1421 | _T_1430; // @[Reg.scala 28:19]
  wire  _T_1433 = _T_1416 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_1434 = _T_1415 & _T_1433; // @[Cache.scala 827:89]
  wire  _T_1435 = _T_1434 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_148 = _T_1435 | _T_1444; // @[Reg.scala 28:19]
  wire  _T_1447 = _T_1416 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_1448 = _T_1415 & _T_1447; // @[Cache.scala 827:89]
  wire  _T_1449 = _T_1448 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_150 = _T_1449 | _T_1458; // @[Reg.scala 28:19]
  wire  _T_1461 = _T_1416 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_1462 = _T_1415 & _T_1461; // @[Cache.scala 827:89]
  wire  _T_1463 = _T_1462 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_152 = _T_1463 | _T_1472; // @[Reg.scala 28:19]
  wire [1:0] _T_1474 = _T_1477 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_1476 = io_cacheOut_r_last_i & _T_189; // @[Cache.scala 824:30]
  wire  _T_1480 = _T_1477 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_1481 = _T_1476 & _T_1480; // @[Cache.scala 827:89]
  wire  _T_1482 = _T_1481 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_155 = _T_1482 | _T_1491; // @[Reg.scala 28:19]
  wire  _T_1494 = _T_1477 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_1495 = _T_1476 & _T_1494; // @[Cache.scala 827:89]
  wire  _T_1496 = _T_1495 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_157 = _T_1496 | _T_1505; // @[Reg.scala 28:19]
  wire  _T_1508 = _T_1477 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_1509 = _T_1476 & _T_1508; // @[Cache.scala 827:89]
  wire  _T_1510 = _T_1509 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_159 = _T_1510 | _T_1519; // @[Reg.scala 28:19]
  wire  _T_1522 = _T_1477 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_1523 = _T_1476 & _T_1522; // @[Cache.scala 827:89]
  wire  _T_1524 = _T_1523 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_161 = _T_1524 | _T_1533; // @[Reg.scala 28:19]
  wire [1:0] _T_1535 = _T_1538 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_1537 = io_cacheOut_r_last_i & _T_191; // @[Cache.scala 824:30]
  wire  _T_1541 = _T_1538 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_1542 = _T_1537 & _T_1541; // @[Cache.scala 827:89]
  wire  _T_1543 = _T_1542 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_164 = _T_1543 | _T_1552; // @[Reg.scala 28:19]
  wire  _T_1555 = _T_1538 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_1556 = _T_1537 & _T_1555; // @[Cache.scala 827:89]
  wire  _T_1557 = _T_1556 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_166 = _T_1557 | _T_1566; // @[Reg.scala 28:19]
  wire  _T_1569 = _T_1538 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_1570 = _T_1537 & _T_1569; // @[Cache.scala 827:89]
  wire  _T_1571 = _T_1570 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_168 = _T_1571 | _T_1580; // @[Reg.scala 28:19]
  wire  _T_1583 = _T_1538 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_1584 = _T_1537 & _T_1583; // @[Cache.scala 827:89]
  wire  _T_1585 = _T_1584 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_170 = _T_1585 | _T_1594; // @[Reg.scala 28:19]
  wire [1:0] _T_1596 = _T_1599 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_1598 = io_cacheOut_r_last_i & _T_193; // @[Cache.scala 824:30]
  wire  _T_1602 = _T_1599 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_1603 = _T_1598 & _T_1602; // @[Cache.scala 827:89]
  wire  _T_1604 = _T_1603 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_173 = _T_1604 | _T_1613; // @[Reg.scala 28:19]
  wire  _T_1616 = _T_1599 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_1617 = _T_1598 & _T_1616; // @[Cache.scala 827:89]
  wire  _T_1618 = _T_1617 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_175 = _T_1618 | _T_1627; // @[Reg.scala 28:19]
  wire  _T_1630 = _T_1599 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_1631 = _T_1598 & _T_1630; // @[Cache.scala 827:89]
  wire  _T_1632 = _T_1631 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_177 = _T_1632 | _T_1641; // @[Reg.scala 28:19]
  wire  _T_1644 = _T_1599 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_1645 = _T_1598 & _T_1644; // @[Cache.scala 827:89]
  wire  _T_1646 = _T_1645 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_179 = _T_1646 | _T_1655; // @[Reg.scala 28:19]
  wire [1:0] _T_1657 = _T_1660 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_1659 = io_cacheOut_r_last_i & _T_195; // @[Cache.scala 824:30]
  wire  _T_1663 = _T_1660 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_1664 = _T_1659 & _T_1663; // @[Cache.scala 827:89]
  wire  _T_1665 = _T_1664 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_182 = _T_1665 | _T_1674; // @[Reg.scala 28:19]
  wire  _T_1677 = _T_1660 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_1678 = _T_1659 & _T_1677; // @[Cache.scala 827:89]
  wire  _T_1679 = _T_1678 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_184 = _T_1679 | _T_1688; // @[Reg.scala 28:19]
  wire  _T_1691 = _T_1660 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_1692 = _T_1659 & _T_1691; // @[Cache.scala 827:89]
  wire  _T_1693 = _T_1692 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_186 = _T_1693 | _T_1702; // @[Reg.scala 28:19]
  wire  _T_1705 = _T_1660 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_1706 = _T_1659 & _T_1705; // @[Cache.scala 827:89]
  wire  _T_1707 = _T_1706 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_188 = _T_1707 | _T_1716; // @[Reg.scala 28:19]
  wire [1:0] _T_1718 = _T_1721 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_1720 = io_cacheOut_r_last_i & _T_197; // @[Cache.scala 824:30]
  wire  _T_1724 = _T_1721 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_1725 = _T_1720 & _T_1724; // @[Cache.scala 827:89]
  wire  _T_1726 = _T_1725 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_191 = _T_1726 | _T_1735; // @[Reg.scala 28:19]
  wire  _T_1738 = _T_1721 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_1739 = _T_1720 & _T_1738; // @[Cache.scala 827:89]
  wire  _T_1740 = _T_1739 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_193 = _T_1740 | _T_1749; // @[Reg.scala 28:19]
  wire  _T_1752 = _T_1721 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_1753 = _T_1720 & _T_1752; // @[Cache.scala 827:89]
  wire  _T_1754 = _T_1753 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_195 = _T_1754 | _T_1763; // @[Reg.scala 28:19]
  wire  _T_1766 = _T_1721 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_1767 = _T_1720 & _T_1766; // @[Cache.scala 827:89]
  wire  _T_1768 = _T_1767 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_197 = _T_1768 | _T_1777; // @[Reg.scala 28:19]
  wire [1:0] _T_1779 = _T_1782 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_1781 = io_cacheOut_r_last_i & _T_199; // @[Cache.scala 824:30]
  wire  _T_1785 = _T_1782 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_1786 = _T_1781 & _T_1785; // @[Cache.scala 827:89]
  wire  _T_1787 = _T_1786 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_200 = _T_1787 | _T_1796; // @[Reg.scala 28:19]
  wire  _T_1799 = _T_1782 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_1800 = _T_1781 & _T_1799; // @[Cache.scala 827:89]
  wire  _T_1801 = _T_1800 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_202 = _T_1801 | _T_1810; // @[Reg.scala 28:19]
  wire  _T_1813 = _T_1782 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_1814 = _T_1781 & _T_1813; // @[Cache.scala 827:89]
  wire  _T_1815 = _T_1814 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_204 = _T_1815 | _T_1824; // @[Reg.scala 28:19]
  wire  _T_1827 = _T_1782 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_1828 = _T_1781 & _T_1827; // @[Cache.scala 827:89]
  wire  _T_1829 = _T_1828 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_206 = _T_1829 | _T_1838; // @[Reg.scala 28:19]
  wire [1:0] _T_1840 = _T_1843 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_1842 = io_cacheOut_r_last_i & _T_201; // @[Cache.scala 824:30]
  wire  _T_1846 = _T_1843 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_1847 = _T_1842 & _T_1846; // @[Cache.scala 827:89]
  wire  _T_1848 = _T_1847 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_209 = _T_1848 | _T_1857; // @[Reg.scala 28:19]
  wire  _T_1860 = _T_1843 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_1861 = _T_1842 & _T_1860; // @[Cache.scala 827:89]
  wire  _T_1862 = _T_1861 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_211 = _T_1862 | _T_1871; // @[Reg.scala 28:19]
  wire  _T_1874 = _T_1843 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_1875 = _T_1842 & _T_1874; // @[Cache.scala 827:89]
  wire  _T_1876 = _T_1875 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_213 = _T_1876 | _T_1885; // @[Reg.scala 28:19]
  wire  _T_1888 = _T_1843 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_1889 = _T_1842 & _T_1888; // @[Cache.scala 827:89]
  wire  _T_1890 = _T_1889 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_215 = _T_1890 | _T_1899; // @[Reg.scala 28:19]
  wire [1:0] _T_1901 = _T_1904 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_1903 = io_cacheOut_r_last_i & _T_203; // @[Cache.scala 824:30]
  wire  _T_1907 = _T_1904 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_1908 = _T_1903 & _T_1907; // @[Cache.scala 827:89]
  wire  _T_1909 = _T_1908 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_218 = _T_1909 | _T_1918; // @[Reg.scala 28:19]
  wire  _T_1921 = _T_1904 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_1922 = _T_1903 & _T_1921; // @[Cache.scala 827:89]
  wire  _T_1923 = _T_1922 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_220 = _T_1923 | _T_1932; // @[Reg.scala 28:19]
  wire  _T_1935 = _T_1904 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_1936 = _T_1903 & _T_1935; // @[Cache.scala 827:89]
  wire  _T_1937 = _T_1936 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_222 = _T_1937 | _T_1946; // @[Reg.scala 28:19]
  wire  _T_1949 = _T_1904 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_1950 = _T_1903 & _T_1949; // @[Cache.scala 827:89]
  wire  _T_1951 = _T_1950 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_224 = _T_1951 | _T_1960; // @[Reg.scala 28:19]
  wire [1:0] _T_1962 = _T_1965 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_1964 = io_cacheOut_r_last_i & _T_205; // @[Cache.scala 824:30]
  wire  _T_1968 = _T_1965 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_1969 = _T_1964 & _T_1968; // @[Cache.scala 827:89]
  wire  _T_1970 = _T_1969 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_227 = _T_1970 | _T_1979; // @[Reg.scala 28:19]
  wire  _T_1982 = _T_1965 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_1983 = _T_1964 & _T_1982; // @[Cache.scala 827:89]
  wire  _T_1984 = _T_1983 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_229 = _T_1984 | _T_1993; // @[Reg.scala 28:19]
  wire  _T_1996 = _T_1965 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_1997 = _T_1964 & _T_1996; // @[Cache.scala 827:89]
  wire  _T_1998 = _T_1997 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_231 = _T_1998 | _T_2007; // @[Reg.scala 28:19]
  wire  _T_2010 = _T_1965 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_2011 = _T_1964 & _T_2010; // @[Cache.scala 827:89]
  wire  _T_2012 = _T_2011 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_233 = _T_2012 | _T_2021; // @[Reg.scala 28:19]
  wire [1:0] _T_2023 = _T_2026 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_2025 = io_cacheOut_r_last_i & _T_207; // @[Cache.scala 824:30]
  wire  _T_2029 = _T_2026 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_2030 = _T_2025 & _T_2029; // @[Cache.scala 827:89]
  wire  _T_2031 = _T_2030 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_236 = _T_2031 | _T_2040; // @[Reg.scala 28:19]
  wire  _T_2043 = _T_2026 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_2044 = _T_2025 & _T_2043; // @[Cache.scala 827:89]
  wire  _T_2045 = _T_2044 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_238 = _T_2045 | _T_2054; // @[Reg.scala 28:19]
  wire  _T_2057 = _T_2026 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_2058 = _T_2025 & _T_2057; // @[Cache.scala 827:89]
  wire  _T_2059 = _T_2058 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_240 = _T_2059 | _T_2068; // @[Reg.scala 28:19]
  wire  _T_2071 = _T_2026 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_2072 = _T_2025 & _T_2071; // @[Cache.scala 827:89]
  wire  _T_2073 = _T_2072 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_242 = _T_2073 | _T_2082; // @[Reg.scala 28:19]
  wire [1:0] _T_2084 = _T_2087 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_2086 = io_cacheOut_r_last_i & _T_209; // @[Cache.scala 824:30]
  wire  _T_2090 = _T_2087 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_2091 = _T_2086 & _T_2090; // @[Cache.scala 827:89]
  wire  _T_2092 = _T_2091 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_245 = _T_2092 | _T_2101; // @[Reg.scala 28:19]
  wire  _T_2104 = _T_2087 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_2105 = _T_2086 & _T_2104; // @[Cache.scala 827:89]
  wire  _T_2106 = _T_2105 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_247 = _T_2106 | _T_2115; // @[Reg.scala 28:19]
  wire  _T_2118 = _T_2087 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_2119 = _T_2086 & _T_2118; // @[Cache.scala 827:89]
  wire  _T_2120 = _T_2119 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_249 = _T_2120 | _T_2129; // @[Reg.scala 28:19]
  wire  _T_2132 = _T_2087 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_2133 = _T_2086 & _T_2132; // @[Cache.scala 827:89]
  wire  _T_2134 = _T_2133 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_251 = _T_2134 | _T_2143; // @[Reg.scala 28:19]
  wire [1:0] _T_2145 = _T_2148 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_2147 = io_cacheOut_r_last_i & _T_211; // @[Cache.scala 824:30]
  wire  _T_2151 = _T_2148 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_2152 = _T_2147 & _T_2151; // @[Cache.scala 827:89]
  wire  _T_2153 = _T_2152 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_254 = _T_2153 | _T_2162; // @[Reg.scala 28:19]
  wire  _T_2165 = _T_2148 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_2166 = _T_2147 & _T_2165; // @[Cache.scala 827:89]
  wire  _T_2167 = _T_2166 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_256 = _T_2167 | _T_2176; // @[Reg.scala 28:19]
  wire  _T_2179 = _T_2148 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_2180 = _T_2147 & _T_2179; // @[Cache.scala 827:89]
  wire  _T_2181 = _T_2180 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_258 = _T_2181 | _T_2190; // @[Reg.scala 28:19]
  wire  _T_2193 = _T_2148 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_2194 = _T_2147 & _T_2193; // @[Cache.scala 827:89]
  wire  _T_2195 = _T_2194 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_260 = _T_2195 | _T_2204; // @[Reg.scala 28:19]
  wire [1:0] _T_2206 = _T_2209 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_2208 = io_cacheOut_r_last_i & _T_213; // @[Cache.scala 824:30]
  wire  _T_2212 = _T_2209 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_2213 = _T_2208 & _T_2212; // @[Cache.scala 827:89]
  wire  _T_2214 = _T_2213 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_263 = _T_2214 | _T_2223; // @[Reg.scala 28:19]
  wire  _T_2226 = _T_2209 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_2227 = _T_2208 & _T_2226; // @[Cache.scala 827:89]
  wire  _T_2228 = _T_2227 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_265 = _T_2228 | _T_2237; // @[Reg.scala 28:19]
  wire  _T_2240 = _T_2209 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_2241 = _T_2208 & _T_2240; // @[Cache.scala 827:89]
  wire  _T_2242 = _T_2241 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_267 = _T_2242 | _T_2251; // @[Reg.scala 28:19]
  wire  _T_2254 = _T_2209 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_2255 = _T_2208 & _T_2254; // @[Cache.scala 827:89]
  wire  _T_2256 = _T_2255 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_269 = _T_2256 | _T_2265; // @[Reg.scala 28:19]
  wire [1:0] _T_2267 = _T_2270 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_2269 = io_cacheOut_r_last_i & _T_215; // @[Cache.scala 824:30]
  wire  _T_2273 = _T_2270 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_2274 = _T_2269 & _T_2273; // @[Cache.scala 827:89]
  wire  _T_2275 = _T_2274 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_272 = _T_2275 | _T_2284; // @[Reg.scala 28:19]
  wire  _T_2287 = _T_2270 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_2288 = _T_2269 & _T_2287; // @[Cache.scala 827:89]
  wire  _T_2289 = _T_2288 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_274 = _T_2289 | _T_2298; // @[Reg.scala 28:19]
  wire  _T_2301 = _T_2270 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_2302 = _T_2269 & _T_2301; // @[Cache.scala 827:89]
  wire  _T_2303 = _T_2302 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_276 = _T_2303 | _T_2312; // @[Reg.scala 28:19]
  wire  _T_2315 = _T_2270 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_2316 = _T_2269 & _T_2315; // @[Cache.scala 827:89]
  wire  _T_2317 = _T_2316 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_278 = _T_2317 | _T_2326; // @[Reg.scala 28:19]
  wire [1:0] _T_2328 = _T_2331 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_2330 = io_cacheOut_r_last_i & _T_217; // @[Cache.scala 824:30]
  wire  _T_2334 = _T_2331 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_2335 = _T_2330 & _T_2334; // @[Cache.scala 827:89]
  wire  _T_2336 = _T_2335 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_281 = _T_2336 | _T_2345; // @[Reg.scala 28:19]
  wire  _T_2348 = _T_2331 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_2349 = _T_2330 & _T_2348; // @[Cache.scala 827:89]
  wire  _T_2350 = _T_2349 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_283 = _T_2350 | _T_2359; // @[Reg.scala 28:19]
  wire  _T_2362 = _T_2331 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_2363 = _T_2330 & _T_2362; // @[Cache.scala 827:89]
  wire  _T_2364 = _T_2363 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_285 = _T_2364 | _T_2373; // @[Reg.scala 28:19]
  wire  _T_2376 = _T_2331 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_2377 = _T_2330 & _T_2376; // @[Cache.scala 827:89]
  wire  _T_2378 = _T_2377 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_287 = _T_2378 | _T_2387; // @[Reg.scala 28:19]
  wire [1:0] _T_2389 = _T_2392 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_2391 = io_cacheOut_r_last_i & _T_219; // @[Cache.scala 824:30]
  wire  _T_2395 = _T_2392 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_2396 = _T_2391 & _T_2395; // @[Cache.scala 827:89]
  wire  _T_2397 = _T_2396 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_290 = _T_2397 | _T_2406; // @[Reg.scala 28:19]
  wire  _T_2409 = _T_2392 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_2410 = _T_2391 & _T_2409; // @[Cache.scala 827:89]
  wire  _T_2411 = _T_2410 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_292 = _T_2411 | _T_2420; // @[Reg.scala 28:19]
  wire  _T_2423 = _T_2392 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_2424 = _T_2391 & _T_2423; // @[Cache.scala 827:89]
  wire  _T_2425 = _T_2424 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_294 = _T_2425 | _T_2434; // @[Reg.scala 28:19]
  wire  _T_2437 = _T_2392 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_2438 = _T_2391 & _T_2437; // @[Cache.scala 827:89]
  wire  _T_2439 = _T_2438 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_296 = _T_2439 | _T_2448; // @[Reg.scala 28:19]
  wire [1:0] _T_2450 = _T_2453 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_2452 = io_cacheOut_r_last_i & _T_221; // @[Cache.scala 824:30]
  wire  _T_2456 = _T_2453 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_2457 = _T_2452 & _T_2456; // @[Cache.scala 827:89]
  wire  _T_2458 = _T_2457 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_299 = _T_2458 | _T_2467; // @[Reg.scala 28:19]
  wire  _T_2470 = _T_2453 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_2471 = _T_2452 & _T_2470; // @[Cache.scala 827:89]
  wire  _T_2472 = _T_2471 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_301 = _T_2472 | _T_2481; // @[Reg.scala 28:19]
  wire  _T_2484 = _T_2453 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_2485 = _T_2452 & _T_2484; // @[Cache.scala 827:89]
  wire  _T_2486 = _T_2485 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_303 = _T_2486 | _T_2495; // @[Reg.scala 28:19]
  wire  _T_2498 = _T_2453 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_2499 = _T_2452 & _T_2498; // @[Cache.scala 827:89]
  wire  _T_2500 = _T_2499 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_305 = _T_2500 | _T_2509; // @[Reg.scala 28:19]
  wire [1:0] _T_2511 = _T_2514 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_2513 = io_cacheOut_r_last_i & _T_223; // @[Cache.scala 824:30]
  wire  _T_2517 = _T_2514 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_2518 = _T_2513 & _T_2517; // @[Cache.scala 827:89]
  wire  _T_2519 = _T_2518 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_308 = _T_2519 | _T_2528; // @[Reg.scala 28:19]
  wire  _T_2531 = _T_2514 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_2532 = _T_2513 & _T_2531; // @[Cache.scala 827:89]
  wire  _T_2533 = _T_2532 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_310 = _T_2533 | _T_2542; // @[Reg.scala 28:19]
  wire  _T_2545 = _T_2514 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_2546 = _T_2513 & _T_2545; // @[Cache.scala 827:89]
  wire  _T_2547 = _T_2546 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_312 = _T_2547 | _T_2556; // @[Reg.scala 28:19]
  wire  _T_2559 = _T_2514 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_2560 = _T_2513 & _T_2559; // @[Cache.scala 827:89]
  wire  _T_2561 = _T_2560 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_314 = _T_2561 | _T_2570; // @[Reg.scala 28:19]
  wire [1:0] _T_2572 = _T_2575 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_2574 = io_cacheOut_r_last_i & _T_225; // @[Cache.scala 824:30]
  wire  _T_2578 = _T_2575 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_2579 = _T_2574 & _T_2578; // @[Cache.scala 827:89]
  wire  _T_2580 = _T_2579 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_317 = _T_2580 | _T_2589; // @[Reg.scala 28:19]
  wire  _T_2592 = _T_2575 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_2593 = _T_2574 & _T_2592; // @[Cache.scala 827:89]
  wire  _T_2594 = _T_2593 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_319 = _T_2594 | _T_2603; // @[Reg.scala 28:19]
  wire  _T_2606 = _T_2575 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_2607 = _T_2574 & _T_2606; // @[Cache.scala 827:89]
  wire  _T_2608 = _T_2607 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_321 = _T_2608 | _T_2617; // @[Reg.scala 28:19]
  wire  _T_2620 = _T_2575 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_2621 = _T_2574 & _T_2620; // @[Cache.scala 827:89]
  wire  _T_2622 = _T_2621 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_323 = _T_2622 | _T_2631; // @[Reg.scala 28:19]
  wire [1:0] _T_2633 = _T_2636 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_2635 = io_cacheOut_r_last_i & _T_227; // @[Cache.scala 824:30]
  wire  _T_2639 = _T_2636 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_2640 = _T_2635 & _T_2639; // @[Cache.scala 827:89]
  wire  _T_2641 = _T_2640 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_326 = _T_2641 | _T_2650; // @[Reg.scala 28:19]
  wire  _T_2653 = _T_2636 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_2654 = _T_2635 & _T_2653; // @[Cache.scala 827:89]
  wire  _T_2655 = _T_2654 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_328 = _T_2655 | _T_2664; // @[Reg.scala 28:19]
  wire  _T_2667 = _T_2636 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_2668 = _T_2635 & _T_2667; // @[Cache.scala 827:89]
  wire  _T_2669 = _T_2668 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_330 = _T_2669 | _T_2678; // @[Reg.scala 28:19]
  wire  _T_2681 = _T_2636 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_2682 = _T_2635 & _T_2681; // @[Cache.scala 827:89]
  wire  _T_2683 = _T_2682 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_332 = _T_2683 | _T_2692; // @[Reg.scala 28:19]
  wire [1:0] _T_2694 = _T_2697 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_2696 = io_cacheOut_r_last_i & _T_229; // @[Cache.scala 824:30]
  wire  _T_2700 = _T_2697 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_2701 = _T_2696 & _T_2700; // @[Cache.scala 827:89]
  wire  _T_2702 = _T_2701 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_335 = _T_2702 | _T_2711; // @[Reg.scala 28:19]
  wire  _T_2714 = _T_2697 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_2715 = _T_2696 & _T_2714; // @[Cache.scala 827:89]
  wire  _T_2716 = _T_2715 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_337 = _T_2716 | _T_2725; // @[Reg.scala 28:19]
  wire  _T_2728 = _T_2697 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_2729 = _T_2696 & _T_2728; // @[Cache.scala 827:89]
  wire  _T_2730 = _T_2729 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_339 = _T_2730 | _T_2739; // @[Reg.scala 28:19]
  wire  _T_2742 = _T_2697 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_2743 = _T_2696 & _T_2742; // @[Cache.scala 827:89]
  wire  _T_2744 = _T_2743 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_341 = _T_2744 | _T_2753; // @[Reg.scala 28:19]
  wire [1:0] _T_2755 = _T_2758 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_2757 = io_cacheOut_r_last_i & _T_231; // @[Cache.scala 824:30]
  wire  _T_2761 = _T_2758 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_2762 = _T_2757 & _T_2761; // @[Cache.scala 827:89]
  wire  _T_2763 = _T_2762 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_344 = _T_2763 | _T_2772; // @[Reg.scala 28:19]
  wire  _T_2775 = _T_2758 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_2776 = _T_2757 & _T_2775; // @[Cache.scala 827:89]
  wire  _T_2777 = _T_2776 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_346 = _T_2777 | _T_2786; // @[Reg.scala 28:19]
  wire  _T_2789 = _T_2758 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_2790 = _T_2757 & _T_2789; // @[Cache.scala 827:89]
  wire  _T_2791 = _T_2790 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_348 = _T_2791 | _T_2800; // @[Reg.scala 28:19]
  wire  _T_2803 = _T_2758 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_2804 = _T_2757 & _T_2803; // @[Cache.scala 827:89]
  wire  _T_2805 = _T_2804 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_350 = _T_2805 | _T_2814; // @[Reg.scala 28:19]
  wire [1:0] _T_2816 = _T_2819 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_2818 = io_cacheOut_r_last_i & _T_233; // @[Cache.scala 824:30]
  wire  _T_2822 = _T_2819 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_2823 = _T_2818 & _T_2822; // @[Cache.scala 827:89]
  wire  _T_2824 = _T_2823 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_353 = _T_2824 | _T_2833; // @[Reg.scala 28:19]
  wire  _T_2836 = _T_2819 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_2837 = _T_2818 & _T_2836; // @[Cache.scala 827:89]
  wire  _T_2838 = _T_2837 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_355 = _T_2838 | _T_2847; // @[Reg.scala 28:19]
  wire  _T_2850 = _T_2819 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_2851 = _T_2818 & _T_2850; // @[Cache.scala 827:89]
  wire  _T_2852 = _T_2851 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_357 = _T_2852 | _T_2861; // @[Reg.scala 28:19]
  wire  _T_2864 = _T_2819 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_2865 = _T_2818 & _T_2864; // @[Cache.scala 827:89]
  wire  _T_2866 = _T_2865 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_359 = _T_2866 | _T_2875; // @[Reg.scala 28:19]
  wire [1:0] _T_2877 = _T_2880 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_2879 = io_cacheOut_r_last_i & _T_235; // @[Cache.scala 824:30]
  wire  _T_2883 = _T_2880 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_2884 = _T_2879 & _T_2883; // @[Cache.scala 827:89]
  wire  _T_2885 = _T_2884 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_362 = _T_2885 | _T_2894; // @[Reg.scala 28:19]
  wire  _T_2897 = _T_2880 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_2898 = _T_2879 & _T_2897; // @[Cache.scala 827:89]
  wire  _T_2899 = _T_2898 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_364 = _T_2899 | _T_2908; // @[Reg.scala 28:19]
  wire  _T_2911 = _T_2880 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_2912 = _T_2879 & _T_2911; // @[Cache.scala 827:89]
  wire  _T_2913 = _T_2912 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_366 = _T_2913 | _T_2922; // @[Reg.scala 28:19]
  wire  _T_2925 = _T_2880 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_2926 = _T_2879 & _T_2925; // @[Cache.scala 827:89]
  wire  _T_2927 = _T_2926 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_368 = _T_2927 | _T_2936; // @[Reg.scala 28:19]
  wire [1:0] _T_2938 = _T_2941 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_2940 = io_cacheOut_r_last_i & _T_237; // @[Cache.scala 824:30]
  wire  _T_2944 = _T_2941 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_2945 = _T_2940 & _T_2944; // @[Cache.scala 827:89]
  wire  _T_2946 = _T_2945 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_371 = _T_2946 | _T_2955; // @[Reg.scala 28:19]
  wire  _T_2958 = _T_2941 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_2959 = _T_2940 & _T_2958; // @[Cache.scala 827:89]
  wire  _T_2960 = _T_2959 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_373 = _T_2960 | _T_2969; // @[Reg.scala 28:19]
  wire  _T_2972 = _T_2941 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_2973 = _T_2940 & _T_2972; // @[Cache.scala 827:89]
  wire  _T_2974 = _T_2973 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_375 = _T_2974 | _T_2983; // @[Reg.scala 28:19]
  wire  _T_2986 = _T_2941 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_2987 = _T_2940 & _T_2986; // @[Cache.scala 827:89]
  wire  _T_2988 = _T_2987 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_377 = _T_2988 | _T_2997; // @[Reg.scala 28:19]
  wire [1:0] _T_2999 = _T_3002 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_3001 = io_cacheOut_r_last_i & _T_239; // @[Cache.scala 824:30]
  wire  _T_3005 = _T_3002 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_3006 = _T_3001 & _T_3005; // @[Cache.scala 827:89]
  wire  _T_3007 = _T_3006 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_380 = _T_3007 | _T_3016; // @[Reg.scala 28:19]
  wire  _T_3019 = _T_3002 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_3020 = _T_3001 & _T_3019; // @[Cache.scala 827:89]
  wire  _T_3021 = _T_3020 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_382 = _T_3021 | _T_3030; // @[Reg.scala 28:19]
  wire  _T_3033 = _T_3002 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_3034 = _T_3001 & _T_3033; // @[Cache.scala 827:89]
  wire  _T_3035 = _T_3034 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_384 = _T_3035 | _T_3044; // @[Reg.scala 28:19]
  wire  _T_3047 = _T_3002 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_3048 = _T_3001 & _T_3047; // @[Cache.scala 827:89]
  wire  _T_3049 = _T_3048 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_386 = _T_3049 | _T_3058; // @[Reg.scala 28:19]
  wire [1:0] _T_3060 = _T_3063 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_3062 = io_cacheOut_r_last_i & _T_241; // @[Cache.scala 824:30]
  wire  _T_3066 = _T_3063 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_3067 = _T_3062 & _T_3066; // @[Cache.scala 827:89]
  wire  _T_3068 = _T_3067 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_389 = _T_3068 | _T_3077; // @[Reg.scala 28:19]
  wire  _T_3080 = _T_3063 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_3081 = _T_3062 & _T_3080; // @[Cache.scala 827:89]
  wire  _T_3082 = _T_3081 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_391 = _T_3082 | _T_3091; // @[Reg.scala 28:19]
  wire  _T_3094 = _T_3063 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_3095 = _T_3062 & _T_3094; // @[Cache.scala 827:89]
  wire  _T_3096 = _T_3095 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_393 = _T_3096 | _T_3105; // @[Reg.scala 28:19]
  wire  _T_3108 = _T_3063 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_3109 = _T_3062 & _T_3108; // @[Cache.scala 827:89]
  wire  _T_3110 = _T_3109 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_395 = _T_3110 | _T_3119; // @[Reg.scala 28:19]
  wire [1:0] _T_3121 = _T_3124 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_3123 = io_cacheOut_r_last_i & _T_243; // @[Cache.scala 824:30]
  wire  _T_3127 = _T_3124 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_3128 = _T_3123 & _T_3127; // @[Cache.scala 827:89]
  wire  _T_3129 = _T_3128 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_398 = _T_3129 | _T_3138; // @[Reg.scala 28:19]
  wire  _T_3141 = _T_3124 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_3142 = _T_3123 & _T_3141; // @[Cache.scala 827:89]
  wire  _T_3143 = _T_3142 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_400 = _T_3143 | _T_3152; // @[Reg.scala 28:19]
  wire  _T_3155 = _T_3124 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_3156 = _T_3123 & _T_3155; // @[Cache.scala 827:89]
  wire  _T_3157 = _T_3156 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_402 = _T_3157 | _T_3166; // @[Reg.scala 28:19]
  wire  _T_3169 = _T_3124 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_3170 = _T_3123 & _T_3169; // @[Cache.scala 827:89]
  wire  _T_3171 = _T_3170 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_404 = _T_3171 | _T_3180; // @[Reg.scala 28:19]
  wire [1:0] _T_3182 = _T_3185 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_3184 = io_cacheOut_r_last_i & _T_245; // @[Cache.scala 824:30]
  wire  _T_3188 = _T_3185 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_3189 = _T_3184 & _T_3188; // @[Cache.scala 827:89]
  wire  _T_3190 = _T_3189 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_407 = _T_3190 | _T_3199; // @[Reg.scala 28:19]
  wire  _T_3202 = _T_3185 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_3203 = _T_3184 & _T_3202; // @[Cache.scala 827:89]
  wire  _T_3204 = _T_3203 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_409 = _T_3204 | _T_3213; // @[Reg.scala 28:19]
  wire  _T_3216 = _T_3185 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_3217 = _T_3184 & _T_3216; // @[Cache.scala 827:89]
  wire  _T_3218 = _T_3217 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_411 = _T_3218 | _T_3227; // @[Reg.scala 28:19]
  wire  _T_3230 = _T_3185 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_3231 = _T_3184 & _T_3230; // @[Cache.scala 827:89]
  wire  _T_3232 = _T_3231 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_413 = _T_3232 | _T_3241; // @[Reg.scala 28:19]
  wire [1:0] _T_3243 = _T_3246 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_3245 = io_cacheOut_r_last_i & _T_247; // @[Cache.scala 824:30]
  wire  _T_3249 = _T_3246 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_3250 = _T_3245 & _T_3249; // @[Cache.scala 827:89]
  wire  _T_3251 = _T_3250 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_416 = _T_3251 | _T_3260; // @[Reg.scala 28:19]
  wire  _T_3263 = _T_3246 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_3264 = _T_3245 & _T_3263; // @[Cache.scala 827:89]
  wire  _T_3265 = _T_3264 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_418 = _T_3265 | _T_3274; // @[Reg.scala 28:19]
  wire  _T_3277 = _T_3246 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_3278 = _T_3245 & _T_3277; // @[Cache.scala 827:89]
  wire  _T_3279 = _T_3278 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_420 = _T_3279 | _T_3288; // @[Reg.scala 28:19]
  wire  _T_3291 = _T_3246 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_3292 = _T_3245 & _T_3291; // @[Cache.scala 827:89]
  wire  _T_3293 = _T_3292 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_422 = _T_3293 | _T_3302; // @[Reg.scala 28:19]
  wire [1:0] _T_3304 = _T_3307 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_3306 = io_cacheOut_r_last_i & _T_249; // @[Cache.scala 824:30]
  wire  _T_3310 = _T_3307 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_3311 = _T_3306 & _T_3310; // @[Cache.scala 827:89]
  wire  _T_3312 = _T_3311 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_425 = _T_3312 | _T_3321; // @[Reg.scala 28:19]
  wire  _T_3324 = _T_3307 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_3325 = _T_3306 & _T_3324; // @[Cache.scala 827:89]
  wire  _T_3326 = _T_3325 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_427 = _T_3326 | _T_3335; // @[Reg.scala 28:19]
  wire  _T_3338 = _T_3307 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_3339 = _T_3306 & _T_3338; // @[Cache.scala 827:89]
  wire  _T_3340 = _T_3339 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_429 = _T_3340 | _T_3349; // @[Reg.scala 28:19]
  wire  _T_3352 = _T_3307 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_3353 = _T_3306 & _T_3352; // @[Cache.scala 827:89]
  wire  _T_3354 = _T_3353 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_431 = _T_3354 | _T_3363; // @[Reg.scala 28:19]
  wire [1:0] _T_3365 = _T_3368 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_3367 = io_cacheOut_r_last_i & _T_251; // @[Cache.scala 824:30]
  wire  _T_3371 = _T_3368 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_3372 = _T_3367 & _T_3371; // @[Cache.scala 827:89]
  wire  _T_3373 = _T_3372 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_434 = _T_3373 | _T_3382; // @[Reg.scala 28:19]
  wire  _T_3385 = _T_3368 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_3386 = _T_3367 & _T_3385; // @[Cache.scala 827:89]
  wire  _T_3387 = _T_3386 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_436 = _T_3387 | _T_3396; // @[Reg.scala 28:19]
  wire  _T_3399 = _T_3368 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_3400 = _T_3367 & _T_3399; // @[Cache.scala 827:89]
  wire  _T_3401 = _T_3400 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_438 = _T_3401 | _T_3410; // @[Reg.scala 28:19]
  wire  _T_3413 = _T_3368 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_3414 = _T_3367 & _T_3413; // @[Cache.scala 827:89]
  wire  _T_3415 = _T_3414 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_440 = _T_3415 | _T_3424; // @[Reg.scala 28:19]
  wire [1:0] _T_3426 = _T_3429 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_3428 = io_cacheOut_r_last_i & _T_253; // @[Cache.scala 824:30]
  wire  _T_3432 = _T_3429 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_3433 = _T_3428 & _T_3432; // @[Cache.scala 827:89]
  wire  _T_3434 = _T_3433 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_443 = _T_3434 | _T_3443; // @[Reg.scala 28:19]
  wire  _T_3446 = _T_3429 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_3447 = _T_3428 & _T_3446; // @[Cache.scala 827:89]
  wire  _T_3448 = _T_3447 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_445 = _T_3448 | _T_3457; // @[Reg.scala 28:19]
  wire  _T_3460 = _T_3429 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_3461 = _T_3428 & _T_3460; // @[Cache.scala 827:89]
  wire  _T_3462 = _T_3461 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_447 = _T_3462 | _T_3471; // @[Reg.scala 28:19]
  wire  _T_3474 = _T_3429 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_3475 = _T_3428 & _T_3474; // @[Cache.scala 827:89]
  wire  _T_3476 = _T_3475 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_449 = _T_3476 | _T_3485; // @[Reg.scala 28:19]
  wire [1:0] _T_3487 = _T_3490 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_3489 = io_cacheOut_r_last_i & _T_255; // @[Cache.scala 824:30]
  wire  _T_3493 = _T_3490 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_3494 = _T_3489 & _T_3493; // @[Cache.scala 827:89]
  wire  _T_3495 = _T_3494 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_452 = _T_3495 | _T_3504; // @[Reg.scala 28:19]
  wire  _T_3507 = _T_3490 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_3508 = _T_3489 & _T_3507; // @[Cache.scala 827:89]
  wire  _T_3509 = _T_3508 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_454 = _T_3509 | _T_3518; // @[Reg.scala 28:19]
  wire  _T_3521 = _T_3490 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_3522 = _T_3489 & _T_3521; // @[Cache.scala 827:89]
  wire  _T_3523 = _T_3522 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_456 = _T_3523 | _T_3532; // @[Reg.scala 28:19]
  wire  _T_3535 = _T_3490 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_3536 = _T_3489 & _T_3535; // @[Cache.scala 827:89]
  wire  _T_3537 = _T_3536 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_458 = _T_3537 | _T_3546; // @[Reg.scala 28:19]
  wire [1:0] _T_3548 = _T_3551 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_3550 = io_cacheOut_r_last_i & _T_257; // @[Cache.scala 824:30]
  wire  _T_3554 = _T_3551 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_3555 = _T_3550 & _T_3554; // @[Cache.scala 827:89]
  wire  _T_3556 = _T_3555 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_461 = _T_3556 | _T_3565; // @[Reg.scala 28:19]
  wire  _T_3568 = _T_3551 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_3569 = _T_3550 & _T_3568; // @[Cache.scala 827:89]
  wire  _T_3570 = _T_3569 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_463 = _T_3570 | _T_3579; // @[Reg.scala 28:19]
  wire  _T_3582 = _T_3551 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_3583 = _T_3550 & _T_3582; // @[Cache.scala 827:89]
  wire  _T_3584 = _T_3583 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_465 = _T_3584 | _T_3593; // @[Reg.scala 28:19]
  wire  _T_3596 = _T_3551 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_3597 = _T_3550 & _T_3596; // @[Cache.scala 827:89]
  wire  _T_3598 = _T_3597 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_467 = _T_3598 | _T_3607; // @[Reg.scala 28:19]
  wire [1:0] _T_3609 = _T_3612 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_3611 = io_cacheOut_r_last_i & _T_259; // @[Cache.scala 824:30]
  wire  _T_3615 = _T_3612 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_3616 = _T_3611 & _T_3615; // @[Cache.scala 827:89]
  wire  _T_3617 = _T_3616 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_470 = _T_3617 | _T_3626; // @[Reg.scala 28:19]
  wire  _T_3629 = _T_3612 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_3630 = _T_3611 & _T_3629; // @[Cache.scala 827:89]
  wire  _T_3631 = _T_3630 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_472 = _T_3631 | _T_3640; // @[Reg.scala 28:19]
  wire  _T_3643 = _T_3612 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_3644 = _T_3611 & _T_3643; // @[Cache.scala 827:89]
  wire  _T_3645 = _T_3644 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_474 = _T_3645 | _T_3654; // @[Reg.scala 28:19]
  wire  _T_3657 = _T_3612 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_3658 = _T_3611 & _T_3657; // @[Cache.scala 827:89]
  wire  _T_3659 = _T_3658 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_476 = _T_3659 | _T_3668; // @[Reg.scala 28:19]
  wire [1:0] _T_3670 = _T_3673 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_3672 = io_cacheOut_r_last_i & _T_261; // @[Cache.scala 824:30]
  wire  _T_3676 = _T_3673 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_3677 = _T_3672 & _T_3676; // @[Cache.scala 827:89]
  wire  _T_3678 = _T_3677 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_479 = _T_3678 | _T_3687; // @[Reg.scala 28:19]
  wire  _T_3690 = _T_3673 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_3691 = _T_3672 & _T_3690; // @[Cache.scala 827:89]
  wire  _T_3692 = _T_3691 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_481 = _T_3692 | _T_3701; // @[Reg.scala 28:19]
  wire  _T_3704 = _T_3673 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_3705 = _T_3672 & _T_3704; // @[Cache.scala 827:89]
  wire  _T_3706 = _T_3705 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_483 = _T_3706 | _T_3715; // @[Reg.scala 28:19]
  wire  _T_3718 = _T_3673 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_3719 = _T_3672 & _T_3718; // @[Cache.scala 827:89]
  wire  _T_3720 = _T_3719 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_485 = _T_3720 | _T_3729; // @[Reg.scala 28:19]
  wire [1:0] _T_3731 = _T_3734 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_3733 = io_cacheOut_r_last_i & _T_263; // @[Cache.scala 824:30]
  wire  _T_3737 = _T_3734 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_3738 = _T_3733 & _T_3737; // @[Cache.scala 827:89]
  wire  _T_3739 = _T_3738 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_488 = _T_3739 | _T_3748; // @[Reg.scala 28:19]
  wire  _T_3751 = _T_3734 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_3752 = _T_3733 & _T_3751; // @[Cache.scala 827:89]
  wire  _T_3753 = _T_3752 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_490 = _T_3753 | _T_3762; // @[Reg.scala 28:19]
  wire  _T_3765 = _T_3734 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_3766 = _T_3733 & _T_3765; // @[Cache.scala 827:89]
  wire  _T_3767 = _T_3766 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_492 = _T_3767 | _T_3776; // @[Reg.scala 28:19]
  wire  _T_3779 = _T_3734 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_3780 = _T_3733 & _T_3779; // @[Cache.scala 827:89]
  wire  _T_3781 = _T_3780 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_494 = _T_3781 | _T_3790; // @[Reg.scala 28:19]
  wire [1:0] _T_3792 = _T_3795 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_3794 = io_cacheOut_r_last_i & _T_265; // @[Cache.scala 824:30]
  wire  _T_3798 = _T_3795 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_3799 = _T_3794 & _T_3798; // @[Cache.scala 827:89]
  wire  _T_3800 = _T_3799 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_497 = _T_3800 | _T_3809; // @[Reg.scala 28:19]
  wire  _T_3812 = _T_3795 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_3813 = _T_3794 & _T_3812; // @[Cache.scala 827:89]
  wire  _T_3814 = _T_3813 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_499 = _T_3814 | _T_3823; // @[Reg.scala 28:19]
  wire  _T_3826 = _T_3795 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_3827 = _T_3794 & _T_3826; // @[Cache.scala 827:89]
  wire  _T_3828 = _T_3827 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_501 = _T_3828 | _T_3837; // @[Reg.scala 28:19]
  wire  _T_3840 = _T_3795 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_3841 = _T_3794 & _T_3840; // @[Cache.scala 827:89]
  wire  _T_3842 = _T_3841 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_503 = _T_3842 | _T_3851; // @[Reg.scala 28:19]
  wire [1:0] _T_3853 = _T_3856 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_3855 = io_cacheOut_r_last_i & _T_267; // @[Cache.scala 824:30]
  wire  _T_3859 = _T_3856 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_3860 = _T_3855 & _T_3859; // @[Cache.scala 827:89]
  wire  _T_3861 = _T_3860 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_506 = _T_3861 | _T_3870; // @[Reg.scala 28:19]
  wire  _T_3873 = _T_3856 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_3874 = _T_3855 & _T_3873; // @[Cache.scala 827:89]
  wire  _T_3875 = _T_3874 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_508 = _T_3875 | _T_3884; // @[Reg.scala 28:19]
  wire  _T_3887 = _T_3856 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_3888 = _T_3855 & _T_3887; // @[Cache.scala 827:89]
  wire  _T_3889 = _T_3888 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_510 = _T_3889 | _T_3898; // @[Reg.scala 28:19]
  wire  _T_3901 = _T_3856 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_3902 = _T_3855 & _T_3901; // @[Cache.scala 827:89]
  wire  _T_3903 = _T_3902 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_512 = _T_3903 | _T_3912; // @[Reg.scala 28:19]
  wire [1:0] _T_3914 = _T_3917 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_3916 = io_cacheOut_r_last_i & _T_269; // @[Cache.scala 824:30]
  wire  _T_3920 = _T_3917 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_3921 = _T_3916 & _T_3920; // @[Cache.scala 827:89]
  wire  _T_3922 = _T_3921 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_515 = _T_3922 | _T_3931; // @[Reg.scala 28:19]
  wire  _T_3934 = _T_3917 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_3935 = _T_3916 & _T_3934; // @[Cache.scala 827:89]
  wire  _T_3936 = _T_3935 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_517 = _T_3936 | _T_3945; // @[Reg.scala 28:19]
  wire  _T_3948 = _T_3917 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_3949 = _T_3916 & _T_3948; // @[Cache.scala 827:89]
  wire  _T_3950 = _T_3949 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_519 = _T_3950 | _T_3959; // @[Reg.scala 28:19]
  wire  _T_3962 = _T_3917 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_3963 = _T_3916 & _T_3962; // @[Cache.scala 827:89]
  wire  _T_3964 = _T_3963 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_521 = _T_3964 | _T_3973; // @[Reg.scala 28:19]
  wire [1:0] _T_3975 = _T_3978 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_3977 = io_cacheOut_r_last_i & _T_271; // @[Cache.scala 824:30]
  wire  _T_3981 = _T_3978 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_3982 = _T_3977 & _T_3981; // @[Cache.scala 827:89]
  wire  _T_3983 = _T_3982 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_524 = _T_3983 | _T_3992; // @[Reg.scala 28:19]
  wire  _T_3995 = _T_3978 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_3996 = _T_3977 & _T_3995; // @[Cache.scala 827:89]
  wire  _T_3997 = _T_3996 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_526 = _T_3997 | _T_4006; // @[Reg.scala 28:19]
  wire  _T_4009 = _T_3978 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_4010 = _T_3977 & _T_4009; // @[Cache.scala 827:89]
  wire  _T_4011 = _T_4010 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_528 = _T_4011 | _T_4020; // @[Reg.scala 28:19]
  wire  _T_4023 = _T_3978 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_4024 = _T_3977 & _T_4023; // @[Cache.scala 827:89]
  wire  _T_4025 = _T_4024 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_530 = _T_4025 | _T_4034; // @[Reg.scala 28:19]
  wire [1:0] _T_4036 = _T_4039 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_4038 = io_cacheOut_r_last_i & _T_273; // @[Cache.scala 824:30]
  wire  _T_4042 = _T_4039 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_4043 = _T_4038 & _T_4042; // @[Cache.scala 827:89]
  wire  _T_4044 = _T_4043 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_533 = _T_4044 | _T_4053; // @[Reg.scala 28:19]
  wire  _T_4056 = _T_4039 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_4057 = _T_4038 & _T_4056; // @[Cache.scala 827:89]
  wire  _T_4058 = _T_4057 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_535 = _T_4058 | _T_4067; // @[Reg.scala 28:19]
  wire  _T_4070 = _T_4039 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_4071 = _T_4038 & _T_4070; // @[Cache.scala 827:89]
  wire  _T_4072 = _T_4071 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_537 = _T_4072 | _T_4081; // @[Reg.scala 28:19]
  wire  _T_4084 = _T_4039 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_4085 = _T_4038 & _T_4084; // @[Cache.scala 827:89]
  wire  _T_4086 = _T_4085 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_539 = _T_4086 | _T_4095; // @[Reg.scala 28:19]
  wire [1:0] _T_4097 = _T_4100 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_4099 = io_cacheOut_r_last_i & _T_275; // @[Cache.scala 824:30]
  wire  _T_4103 = _T_4100 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_4104 = _T_4099 & _T_4103; // @[Cache.scala 827:89]
  wire  _T_4105 = _T_4104 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_542 = _T_4105 | _T_4114; // @[Reg.scala 28:19]
  wire  _T_4117 = _T_4100 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_4118 = _T_4099 & _T_4117; // @[Cache.scala 827:89]
  wire  _T_4119 = _T_4118 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_544 = _T_4119 | _T_4128; // @[Reg.scala 28:19]
  wire  _T_4131 = _T_4100 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_4132 = _T_4099 & _T_4131; // @[Cache.scala 827:89]
  wire  _T_4133 = _T_4132 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_546 = _T_4133 | _T_4142; // @[Reg.scala 28:19]
  wire  _T_4145 = _T_4100 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_4146 = _T_4099 & _T_4145; // @[Cache.scala 827:89]
  wire  _T_4147 = _T_4146 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_548 = _T_4147 | _T_4156; // @[Reg.scala 28:19]
  wire [1:0] _T_4158 = _T_4161 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_4160 = io_cacheOut_r_last_i & _T_277; // @[Cache.scala 824:30]
  wire  _T_4164 = _T_4161 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_4165 = _T_4160 & _T_4164; // @[Cache.scala 827:89]
  wire  _T_4166 = _T_4165 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_551 = _T_4166 | _T_4175; // @[Reg.scala 28:19]
  wire  _T_4178 = _T_4161 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_4179 = _T_4160 & _T_4178; // @[Cache.scala 827:89]
  wire  _T_4180 = _T_4179 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_553 = _T_4180 | _T_4189; // @[Reg.scala 28:19]
  wire  _T_4192 = _T_4161 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_4193 = _T_4160 & _T_4192; // @[Cache.scala 827:89]
  wire  _T_4194 = _T_4193 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_555 = _T_4194 | _T_4203; // @[Reg.scala 28:19]
  wire  _T_4206 = _T_4161 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_4207 = _T_4160 & _T_4206; // @[Cache.scala 827:89]
  wire  _T_4208 = _T_4207 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_557 = _T_4208 | _T_4217; // @[Reg.scala 28:19]
  wire [1:0] _T_4219 = _T_4222 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_4221 = io_cacheOut_r_last_i & _T_279; // @[Cache.scala 824:30]
  wire  _T_4225 = _T_4222 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_4226 = _T_4221 & _T_4225; // @[Cache.scala 827:89]
  wire  _T_4227 = _T_4226 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_560 = _T_4227 | _T_4236; // @[Reg.scala 28:19]
  wire  _T_4239 = _T_4222 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_4240 = _T_4221 & _T_4239; // @[Cache.scala 827:89]
  wire  _T_4241 = _T_4240 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_562 = _T_4241 | _T_4250; // @[Reg.scala 28:19]
  wire  _T_4253 = _T_4222 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_4254 = _T_4221 & _T_4253; // @[Cache.scala 827:89]
  wire  _T_4255 = _T_4254 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_564 = _T_4255 | _T_4264; // @[Reg.scala 28:19]
  wire  _T_4267 = _T_4222 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_4268 = _T_4221 & _T_4267; // @[Cache.scala 827:89]
  wire  _T_4269 = _T_4268 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_566 = _T_4269 | _T_4278; // @[Reg.scala 28:19]
  wire [1:0] _T_4280 = _T_4283 + 2'h1; // @[Cache.scala 822:25]
  wire  _T_4282 = io_cacheOut_r_last_i & _T_281; // @[Cache.scala 824:30]
  wire  _T_4286 = _T_4283 == 2'h0; // @[Cache.scala 827:108]
  wire  _T_4287 = _T_4282 & _T_4286; // @[Cache.scala 827:89]
  wire  _T_4288 = _T_4287 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_569 = _T_4288 | _T_4297; // @[Reg.scala 28:19]
  wire  _T_4300 = _T_4283 == 2'h1; // @[Cache.scala 827:108]
  wire  _T_4301 = _T_4282 & _T_4300; // @[Cache.scala 827:89]
  wire  _T_4302 = _T_4301 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_571 = _T_4302 | _T_4311; // @[Reg.scala 28:19]
  wire  _T_4314 = _T_4283 == 2'h2; // @[Cache.scala 827:108]
  wire  _T_4315 = _T_4282 & _T_4314; // @[Cache.scala 827:89]
  wire  _T_4316 = _T_4315 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_573 = _T_4316 | _T_4325; // @[Reg.scala 28:19]
  wire  _T_4328 = _T_4283 == 2'h3; // @[Cache.scala 827:108]
  wire  _T_4329 = _T_4282 & _T_4328; // @[Cache.scala 827:89]
  wire  _T_4330 = _T_4329 & _T_25; // @[Cache.scala 827:116]
  wire  _GEN_575 = _T_4330 | _T_4339; // @[Reg.scala 28:19]
  wire [7:0] _T_4344 = io_cacheIn_mask[0] ? 8'h0 : 8'hff; // @[Cache.scala 840:26]
  wire [7:0] _T_4348 = io_cacheIn_mask[1] ? 8'h0 : 8'hff; // @[Cache.scala 840:26]
  wire [7:0] _T_4352 = io_cacheIn_mask[2] ? 8'h0 : 8'hff; // @[Cache.scala 840:26]
  wire [7:0] _T_4356 = io_cacheIn_mask[3] ? 8'h0 : 8'hff; // @[Cache.scala 840:26]
  wire [7:0] _T_4360 = io_cacheIn_mask[4] ? 8'h0 : 8'hff; // @[Cache.scala 840:26]
  wire [7:0] _T_4364 = io_cacheIn_mask[5] ? 8'h0 : 8'hff; // @[Cache.scala 840:26]
  wire [7:0] _T_4368 = io_cacheIn_mask[6] ? 8'h0 : 8'hff; // @[Cache.scala 840:26]
  wire [7:0] _T_4372 = io_cacheIn_mask[7] ? 8'h0 : 8'hff; // @[Cache.scala 840:26]
  wire [127:0] _T_4383 = {_T_4372,_T_4368,_T_4364,_T_4360,_T_4356,_T_4352,_T_4348,_T_4344,64'hffffffffffffffff}; // @[Cat.scala 29:58]
  wire [127:0] _T_4393 = {64'hffffffffffffffff,_T_4372,_T_4368,_T_4364,_T_4360,_T_4356,_T_4352,_T_4348,_T_4344}; // @[Cat.scala 29:58]
  wire [127:0] _T_4394 = io_cacheIn_addr[3] ? _T_4383 : _T_4393; // @[Cache.scala 847:27]
  wire  _T_4395 = io_cacheIn_valid & io_cacheIn_wen; // @[Cache.scala 865:48]
  wire  _T_4397 = io_cacheIn_valid & _T_284; // @[Cache.scala 875:38]
  wire  _T_4398 = _T_4397 & _T_24; // @[Cache.scala 875:55]
  wire  _T_4399 = _T_25 & io_cacheOut_r_valid_i; // @[Cache.scala 875:78]
  wire  _T_4400 = 2'h0 == _T_433; // @[Cache.scala 875:113]
  wire  _T_4401 = _T_4399 & _T_4400; // @[Cache.scala 875:104]
  wire  _T_4402 = _T_4398 | _T_4401; // @[Cache.scala 875:66]
  wire  _T_4404 = io_cacheIn_wen & _T_24; // @[Cache.scala 877:36]
  wire  _T_4408 = _T_4404 | _T_4401; // @[Cache.scala 877:47]
  wire [127:0] _T_4410 = {io_cacheOut_r_data_i,64'h0}; // @[Cat.scala 29:58]
  wire [127:0] _T_4411 = {64'h0,io_cacheOut_r_data_i}; // @[Cat.scala 29:58]
  wire [127:0] _T_4412 = io_cacheOut_r_last_i ? _T_4410 : _T_4411; // @[Cache.scala 880:12]
  wire [127:0] _T_4414 = {io_cacheIn_data_write,64'h0}; // @[Cat.scala 29:58]
  wire [127:0] _T_4415 = {64'h0,io_cacheIn_data_write}; // @[Cat.scala 29:58]
  wire [127:0] _T_4416 = io_cacheIn_addr[3] ? _T_4414 : _T_4415; // @[Cache.scala 881:12]
  wire [127:0] _T_4424 = io_cacheOut_r_last_i ? 128'hffffffffffffffff : 128'hffffffffffffffff0000000000000000; // @[Cache.scala 885:12]
  wire  _T_4426 = io_cacheIn_valid & _T_286; // @[Cache.scala 875:38]
  wire  _T_4427 = _T_4426 & _T_24; // @[Cache.scala 875:55]
  wire  _T_4429 = 2'h1 == _T_433; // @[Cache.scala 875:113]
  wire  _T_4430 = _T_4399 & _T_4429; // @[Cache.scala 875:104]
  wire  _T_4431 = _T_4427 | _T_4430; // @[Cache.scala 875:66]
  wire  _T_4437 = _T_4404 | _T_4430; // @[Cache.scala 877:47]
  wire  _T_4455 = io_cacheIn_valid & _T_288; // @[Cache.scala 875:38]
  wire  _T_4456 = _T_4455 & _T_24; // @[Cache.scala 875:55]
  wire  _T_4458 = 2'h2 == _T_433; // @[Cache.scala 875:113]
  wire  _T_4459 = _T_4399 & _T_4458; // @[Cache.scala 875:104]
  wire  _T_4460 = _T_4456 | _T_4459; // @[Cache.scala 875:66]
  wire  _T_4466 = _T_4404 | _T_4459; // @[Cache.scala 877:47]
  wire  _T_4484 = io_cacheIn_valid & _T_290; // @[Cache.scala 875:38]
  wire  _T_4485 = _T_4484 & _T_24; // @[Cache.scala 875:55]
  wire  _T_4487 = 2'h3 == _T_433; // @[Cache.scala 875:113]
  wire  _T_4488 = _T_4399 & _T_4487; // @[Cache.scala 875:104]
  wire  _T_4489 = _T_4485 | _T_4488; // @[Cache.scala 875:66]
  wire  _T_4495 = _T_4404 | _T_4488; // @[Cache.scala 877:47]
  wire  _T_4513 = _T_27 & io_cacheOut_w_ready_i; // @[Cache.scala 891:33]
  wire  _T_4514 = _T_4513 | _T_28; // @[Cache.scala 891:58]
  assign io_cacheOut_ar_valid_o = _T_4 == 3'h1; // @[Cache.scala 808:28]
  assign io_cacheOut_ar_addr_o = {io_cacheIn_addr[31:4],4'h0}; // @[Cache.scala 807:27]
  assign io_cacheOut_ar_len_o = {{7'd0}, _T_25}; // @[Cache.scala 806:26]
  assign io_cacheOut_w_valid_o = _T_4395 & _T_24; // @[Cache.scala 865:27]
  assign io_cacheOut_w_data_o = io_cacheIn_data_write; // @[Cache.scala 866:26]
  assign io_cacheOut_w_addr_o = io_cacheIn_addr; // @[Cache.scala 867:26]
  assign io_cacheOut_w_mask_o = io_cacheIn_mask; // @[Cache.scala 868:26]
  assign io_cacheOut_wsize = io_cacheIn_rsize; // @[Cache.scala 893:23]
  assign io_cacheIn_ready = _T_4514 | _T_26; // @[Cache.scala 891:22]
  assign io_cacheIn_data_read = io_cacheIn_addr[3] ? _T_301[127:64] : _T_301[63:0]; // @[Cache.scala 792:26]
  assign io_SRAMIO_0_cen = ~_T_4402; // @[Cache.scala 875:15]
  assign io_SRAMIO_0_wen = ~_T_4408; // @[Cache.scala 877:15]
  assign io_SRAMIO_0_wdata = _T_25 ? _T_4412 : _T_4416; // @[Cache.scala 878:17]
  assign io_SRAMIO_0_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 876:16]
  assign io_SRAMIO_0_wmask = _T_25 ? _T_4424 : _T_4394; // @[Cache.scala 883:17]
  assign io_SRAMIO_1_cen = ~_T_4431; // @[Cache.scala 875:15]
  assign io_SRAMIO_1_wen = ~_T_4437; // @[Cache.scala 877:15]
  assign io_SRAMIO_1_wdata = _T_25 ? _T_4412 : _T_4416; // @[Cache.scala 878:17]
  assign io_SRAMIO_1_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 876:16]
  assign io_SRAMIO_1_wmask = _T_25 ? _T_4424 : _T_4394; // @[Cache.scala 883:17]
  assign io_SRAMIO_2_cen = ~_T_4460; // @[Cache.scala 875:15]
  assign io_SRAMIO_2_wen = ~_T_4466; // @[Cache.scala 877:15]
  assign io_SRAMIO_2_wdata = _T_25 ? _T_4412 : _T_4416; // @[Cache.scala 878:17]
  assign io_SRAMIO_2_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 876:16]
  assign io_SRAMIO_2_wmask = _T_25 ? _T_4424 : _T_4394; // @[Cache.scala 883:17]
  assign io_SRAMIO_3_cen = ~_T_4489; // @[Cache.scala 875:15]
  assign io_SRAMIO_3_wen = ~_T_4495; // @[Cache.scala 877:15]
  assign io_SRAMIO_3_wdata = _T_25 ? _T_4412 : _T_4416; // @[Cache.scala 878:17]
  assign io_SRAMIO_3_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 876:16]
  assign io_SRAMIO_3_wmask = _T_25 ? _T_4424 : _T_4394; // @[Cache.scala 883:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_4 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  _T_4297 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_4236 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _T_4175 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_4114 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_4053 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_3992 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_3931 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_3870 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_3809 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_3748 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_3687 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_3626 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_3565 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_3504 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_3443 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _T_3382 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _T_3321 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_3260 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _T_3199 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _T_3138 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_3077 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  _T_3016 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _T_2955 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  _T_2894 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  _T_2833 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  _T_2772 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  _T_2711 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  _T_2650 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  _T_2589 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  _T_2528 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  _T_2467 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  _T_2406 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  _T_2345 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  _T_2284 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  _T_2223 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  _T_2162 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  _T_2101 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  _T_2040 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  _T_1979 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  _T_1918 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  _T_1857 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  _T_1796 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  _T_1735 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  _T_1674 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  _T_1613 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  _T_1552 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  _T_1491 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  _T_1430 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  _T_1369 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  _T_1308 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  _T_1247 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  _T_1186 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  _T_1125 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  _T_1064 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  _T_1003 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  _T_942 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  _T_881 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  _T_820 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  _T_759 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  _T_698 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  _T_637 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  _T_576 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  _T_515 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  _T_454 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  _T_4289 = _RAND_65[21:0];
  _RAND_66 = {1{`RANDOM}};
  _T_4228 = _RAND_66[21:0];
  _RAND_67 = {1{`RANDOM}};
  _T_4167 = _RAND_67[21:0];
  _RAND_68 = {1{`RANDOM}};
  _T_4106 = _RAND_68[21:0];
  _RAND_69 = {1{`RANDOM}};
  _T_4045 = _RAND_69[21:0];
  _RAND_70 = {1{`RANDOM}};
  _T_3984 = _RAND_70[21:0];
  _RAND_71 = {1{`RANDOM}};
  _T_3923 = _RAND_71[21:0];
  _RAND_72 = {1{`RANDOM}};
  _T_3862 = _RAND_72[21:0];
  _RAND_73 = {1{`RANDOM}};
  _T_3801 = _RAND_73[21:0];
  _RAND_74 = {1{`RANDOM}};
  _T_3740 = _RAND_74[21:0];
  _RAND_75 = {1{`RANDOM}};
  _T_3679 = _RAND_75[21:0];
  _RAND_76 = {1{`RANDOM}};
  _T_3618 = _RAND_76[21:0];
  _RAND_77 = {1{`RANDOM}};
  _T_3557 = _RAND_77[21:0];
  _RAND_78 = {1{`RANDOM}};
  _T_3496 = _RAND_78[21:0];
  _RAND_79 = {1{`RANDOM}};
  _T_3435 = _RAND_79[21:0];
  _RAND_80 = {1{`RANDOM}};
  _T_3374 = _RAND_80[21:0];
  _RAND_81 = {1{`RANDOM}};
  _T_3313 = _RAND_81[21:0];
  _RAND_82 = {1{`RANDOM}};
  _T_3252 = _RAND_82[21:0];
  _RAND_83 = {1{`RANDOM}};
  _T_3191 = _RAND_83[21:0];
  _RAND_84 = {1{`RANDOM}};
  _T_3130 = _RAND_84[21:0];
  _RAND_85 = {1{`RANDOM}};
  _T_3069 = _RAND_85[21:0];
  _RAND_86 = {1{`RANDOM}};
  _T_3008 = _RAND_86[21:0];
  _RAND_87 = {1{`RANDOM}};
  _T_2947 = _RAND_87[21:0];
  _RAND_88 = {1{`RANDOM}};
  _T_2886 = _RAND_88[21:0];
  _RAND_89 = {1{`RANDOM}};
  _T_2825 = _RAND_89[21:0];
  _RAND_90 = {1{`RANDOM}};
  _T_2764 = _RAND_90[21:0];
  _RAND_91 = {1{`RANDOM}};
  _T_2703 = _RAND_91[21:0];
  _RAND_92 = {1{`RANDOM}};
  _T_2642 = _RAND_92[21:0];
  _RAND_93 = {1{`RANDOM}};
  _T_2581 = _RAND_93[21:0];
  _RAND_94 = {1{`RANDOM}};
  _T_2520 = _RAND_94[21:0];
  _RAND_95 = {1{`RANDOM}};
  _T_2459 = _RAND_95[21:0];
  _RAND_96 = {1{`RANDOM}};
  _T_2398 = _RAND_96[21:0];
  _RAND_97 = {1{`RANDOM}};
  _T_2337 = _RAND_97[21:0];
  _RAND_98 = {1{`RANDOM}};
  _T_2276 = _RAND_98[21:0];
  _RAND_99 = {1{`RANDOM}};
  _T_2215 = _RAND_99[21:0];
  _RAND_100 = {1{`RANDOM}};
  _T_2154 = _RAND_100[21:0];
  _RAND_101 = {1{`RANDOM}};
  _T_2093 = _RAND_101[21:0];
  _RAND_102 = {1{`RANDOM}};
  _T_2032 = _RAND_102[21:0];
  _RAND_103 = {1{`RANDOM}};
  _T_1971 = _RAND_103[21:0];
  _RAND_104 = {1{`RANDOM}};
  _T_1910 = _RAND_104[21:0];
  _RAND_105 = {1{`RANDOM}};
  _T_1849 = _RAND_105[21:0];
  _RAND_106 = {1{`RANDOM}};
  _T_1788 = _RAND_106[21:0];
  _RAND_107 = {1{`RANDOM}};
  _T_1727 = _RAND_107[21:0];
  _RAND_108 = {1{`RANDOM}};
  _T_1666 = _RAND_108[21:0];
  _RAND_109 = {1{`RANDOM}};
  _T_1605 = _RAND_109[21:0];
  _RAND_110 = {1{`RANDOM}};
  _T_1544 = _RAND_110[21:0];
  _RAND_111 = {1{`RANDOM}};
  _T_1483 = _RAND_111[21:0];
  _RAND_112 = {1{`RANDOM}};
  _T_1422 = _RAND_112[21:0];
  _RAND_113 = {1{`RANDOM}};
  _T_1361 = _RAND_113[21:0];
  _RAND_114 = {1{`RANDOM}};
  _T_1300 = _RAND_114[21:0];
  _RAND_115 = {1{`RANDOM}};
  _T_1239 = _RAND_115[21:0];
  _RAND_116 = {1{`RANDOM}};
  _T_1178 = _RAND_116[21:0];
  _RAND_117 = {1{`RANDOM}};
  _T_1117 = _RAND_117[21:0];
  _RAND_118 = {1{`RANDOM}};
  _T_1056 = _RAND_118[21:0];
  _RAND_119 = {1{`RANDOM}};
  _T_995 = _RAND_119[21:0];
  _RAND_120 = {1{`RANDOM}};
  _T_934 = _RAND_120[21:0];
  _RAND_121 = {1{`RANDOM}};
  _T_873 = _RAND_121[21:0];
  _RAND_122 = {1{`RANDOM}};
  _T_812 = _RAND_122[21:0];
  _RAND_123 = {1{`RANDOM}};
  _T_751 = _RAND_123[21:0];
  _RAND_124 = {1{`RANDOM}};
  _T_690 = _RAND_124[21:0];
  _RAND_125 = {1{`RANDOM}};
  _T_629 = _RAND_125[21:0];
  _RAND_126 = {1{`RANDOM}};
  _T_568 = _RAND_126[21:0];
  _RAND_127 = {1{`RANDOM}};
  _T_507 = _RAND_127[21:0];
  _RAND_128 = {1{`RANDOM}};
  _T_446 = _RAND_128[21:0];
  _RAND_129 = {1{`RANDOM}};
  _T_4311 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  _T_4250 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  _T_4189 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  _T_4128 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  _T_4067 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  _T_4006 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  _T_3945 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  _T_3884 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  _T_3823 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  _T_3762 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  _T_3701 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  _T_3640 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  _T_3579 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  _T_3518 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  _T_3457 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  _T_3396 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  _T_3335 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  _T_3274 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  _T_3213 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  _T_3152 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  _T_3091 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  _T_3030 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  _T_2969 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  _T_2908 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  _T_2847 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  _T_2786 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  _T_2725 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  _T_2664 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  _T_2603 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  _T_2542 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  _T_2481 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  _T_2420 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  _T_2359 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  _T_2298 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  _T_2237 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  _T_2176 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  _T_2115 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  _T_2054 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  _T_1993 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  _T_1932 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  _T_1871 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  _T_1810 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  _T_1749 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  _T_1688 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  _T_1627 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  _T_1566 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  _T_1505 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  _T_1444 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  _T_1383 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  _T_1322 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  _T_1261 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  _T_1200 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  _T_1139 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  _T_1078 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  _T_1017 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  _T_956 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  _T_895 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  _T_834 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  _T_773 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  _T_712 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  _T_651 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  _T_590 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  _T_529 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  _T_468 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  _T_4303 = _RAND_193[21:0];
  _RAND_194 = {1{`RANDOM}};
  _T_4242 = _RAND_194[21:0];
  _RAND_195 = {1{`RANDOM}};
  _T_4181 = _RAND_195[21:0];
  _RAND_196 = {1{`RANDOM}};
  _T_4120 = _RAND_196[21:0];
  _RAND_197 = {1{`RANDOM}};
  _T_4059 = _RAND_197[21:0];
  _RAND_198 = {1{`RANDOM}};
  _T_3998 = _RAND_198[21:0];
  _RAND_199 = {1{`RANDOM}};
  _T_3937 = _RAND_199[21:0];
  _RAND_200 = {1{`RANDOM}};
  _T_3876 = _RAND_200[21:0];
  _RAND_201 = {1{`RANDOM}};
  _T_3815 = _RAND_201[21:0];
  _RAND_202 = {1{`RANDOM}};
  _T_3754 = _RAND_202[21:0];
  _RAND_203 = {1{`RANDOM}};
  _T_3693 = _RAND_203[21:0];
  _RAND_204 = {1{`RANDOM}};
  _T_3632 = _RAND_204[21:0];
  _RAND_205 = {1{`RANDOM}};
  _T_3571 = _RAND_205[21:0];
  _RAND_206 = {1{`RANDOM}};
  _T_3510 = _RAND_206[21:0];
  _RAND_207 = {1{`RANDOM}};
  _T_3449 = _RAND_207[21:0];
  _RAND_208 = {1{`RANDOM}};
  _T_3388 = _RAND_208[21:0];
  _RAND_209 = {1{`RANDOM}};
  _T_3327 = _RAND_209[21:0];
  _RAND_210 = {1{`RANDOM}};
  _T_3266 = _RAND_210[21:0];
  _RAND_211 = {1{`RANDOM}};
  _T_3205 = _RAND_211[21:0];
  _RAND_212 = {1{`RANDOM}};
  _T_3144 = _RAND_212[21:0];
  _RAND_213 = {1{`RANDOM}};
  _T_3083 = _RAND_213[21:0];
  _RAND_214 = {1{`RANDOM}};
  _T_3022 = _RAND_214[21:0];
  _RAND_215 = {1{`RANDOM}};
  _T_2961 = _RAND_215[21:0];
  _RAND_216 = {1{`RANDOM}};
  _T_2900 = _RAND_216[21:0];
  _RAND_217 = {1{`RANDOM}};
  _T_2839 = _RAND_217[21:0];
  _RAND_218 = {1{`RANDOM}};
  _T_2778 = _RAND_218[21:0];
  _RAND_219 = {1{`RANDOM}};
  _T_2717 = _RAND_219[21:0];
  _RAND_220 = {1{`RANDOM}};
  _T_2656 = _RAND_220[21:0];
  _RAND_221 = {1{`RANDOM}};
  _T_2595 = _RAND_221[21:0];
  _RAND_222 = {1{`RANDOM}};
  _T_2534 = _RAND_222[21:0];
  _RAND_223 = {1{`RANDOM}};
  _T_2473 = _RAND_223[21:0];
  _RAND_224 = {1{`RANDOM}};
  _T_2412 = _RAND_224[21:0];
  _RAND_225 = {1{`RANDOM}};
  _T_2351 = _RAND_225[21:0];
  _RAND_226 = {1{`RANDOM}};
  _T_2290 = _RAND_226[21:0];
  _RAND_227 = {1{`RANDOM}};
  _T_2229 = _RAND_227[21:0];
  _RAND_228 = {1{`RANDOM}};
  _T_2168 = _RAND_228[21:0];
  _RAND_229 = {1{`RANDOM}};
  _T_2107 = _RAND_229[21:0];
  _RAND_230 = {1{`RANDOM}};
  _T_2046 = _RAND_230[21:0];
  _RAND_231 = {1{`RANDOM}};
  _T_1985 = _RAND_231[21:0];
  _RAND_232 = {1{`RANDOM}};
  _T_1924 = _RAND_232[21:0];
  _RAND_233 = {1{`RANDOM}};
  _T_1863 = _RAND_233[21:0];
  _RAND_234 = {1{`RANDOM}};
  _T_1802 = _RAND_234[21:0];
  _RAND_235 = {1{`RANDOM}};
  _T_1741 = _RAND_235[21:0];
  _RAND_236 = {1{`RANDOM}};
  _T_1680 = _RAND_236[21:0];
  _RAND_237 = {1{`RANDOM}};
  _T_1619 = _RAND_237[21:0];
  _RAND_238 = {1{`RANDOM}};
  _T_1558 = _RAND_238[21:0];
  _RAND_239 = {1{`RANDOM}};
  _T_1497 = _RAND_239[21:0];
  _RAND_240 = {1{`RANDOM}};
  _T_1436 = _RAND_240[21:0];
  _RAND_241 = {1{`RANDOM}};
  _T_1375 = _RAND_241[21:0];
  _RAND_242 = {1{`RANDOM}};
  _T_1314 = _RAND_242[21:0];
  _RAND_243 = {1{`RANDOM}};
  _T_1253 = _RAND_243[21:0];
  _RAND_244 = {1{`RANDOM}};
  _T_1192 = _RAND_244[21:0];
  _RAND_245 = {1{`RANDOM}};
  _T_1131 = _RAND_245[21:0];
  _RAND_246 = {1{`RANDOM}};
  _T_1070 = _RAND_246[21:0];
  _RAND_247 = {1{`RANDOM}};
  _T_1009 = _RAND_247[21:0];
  _RAND_248 = {1{`RANDOM}};
  _T_948 = _RAND_248[21:0];
  _RAND_249 = {1{`RANDOM}};
  _T_887 = _RAND_249[21:0];
  _RAND_250 = {1{`RANDOM}};
  _T_826 = _RAND_250[21:0];
  _RAND_251 = {1{`RANDOM}};
  _T_765 = _RAND_251[21:0];
  _RAND_252 = {1{`RANDOM}};
  _T_704 = _RAND_252[21:0];
  _RAND_253 = {1{`RANDOM}};
  _T_643 = _RAND_253[21:0];
  _RAND_254 = {1{`RANDOM}};
  _T_582 = _RAND_254[21:0];
  _RAND_255 = {1{`RANDOM}};
  _T_521 = _RAND_255[21:0];
  _RAND_256 = {1{`RANDOM}};
  _T_460 = _RAND_256[21:0];
  _RAND_257 = {1{`RANDOM}};
  _T_4325 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  _T_4264 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  _T_4203 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  _T_4142 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  _T_4081 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  _T_4020 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  _T_3959 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  _T_3898 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  _T_3837 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  _T_3776 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  _T_3715 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  _T_3654 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  _T_3593 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  _T_3532 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  _T_3471 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  _T_3410 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  _T_3349 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  _T_3288 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  _T_3227 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  _T_3166 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  _T_3105 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  _T_3044 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  _T_2983 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  _T_2922 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  _T_2861 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  _T_2800 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  _T_2739 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  _T_2678 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  _T_2617 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  _T_2556 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  _T_2495 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  _T_2434 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  _T_2373 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  _T_2312 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  _T_2251 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  _T_2190 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  _T_2129 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  _T_2068 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  _T_2007 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  _T_1946 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  _T_1885 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  _T_1824 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  _T_1763 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  _T_1702 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  _T_1641 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  _T_1580 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  _T_1519 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  _T_1458 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  _T_1397 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  _T_1336 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  _T_1275 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  _T_1214 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  _T_1153 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  _T_1092 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  _T_1031 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  _T_970 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  _T_909 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  _T_848 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  _T_787 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  _T_726 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  _T_665 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  _T_604 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  _T_543 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  _T_482 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  _T_4317 = _RAND_321[21:0];
  _RAND_322 = {1{`RANDOM}};
  _T_4256 = _RAND_322[21:0];
  _RAND_323 = {1{`RANDOM}};
  _T_4195 = _RAND_323[21:0];
  _RAND_324 = {1{`RANDOM}};
  _T_4134 = _RAND_324[21:0];
  _RAND_325 = {1{`RANDOM}};
  _T_4073 = _RAND_325[21:0];
  _RAND_326 = {1{`RANDOM}};
  _T_4012 = _RAND_326[21:0];
  _RAND_327 = {1{`RANDOM}};
  _T_3951 = _RAND_327[21:0];
  _RAND_328 = {1{`RANDOM}};
  _T_3890 = _RAND_328[21:0];
  _RAND_329 = {1{`RANDOM}};
  _T_3829 = _RAND_329[21:0];
  _RAND_330 = {1{`RANDOM}};
  _T_3768 = _RAND_330[21:0];
  _RAND_331 = {1{`RANDOM}};
  _T_3707 = _RAND_331[21:0];
  _RAND_332 = {1{`RANDOM}};
  _T_3646 = _RAND_332[21:0];
  _RAND_333 = {1{`RANDOM}};
  _T_3585 = _RAND_333[21:0];
  _RAND_334 = {1{`RANDOM}};
  _T_3524 = _RAND_334[21:0];
  _RAND_335 = {1{`RANDOM}};
  _T_3463 = _RAND_335[21:0];
  _RAND_336 = {1{`RANDOM}};
  _T_3402 = _RAND_336[21:0];
  _RAND_337 = {1{`RANDOM}};
  _T_3341 = _RAND_337[21:0];
  _RAND_338 = {1{`RANDOM}};
  _T_3280 = _RAND_338[21:0];
  _RAND_339 = {1{`RANDOM}};
  _T_3219 = _RAND_339[21:0];
  _RAND_340 = {1{`RANDOM}};
  _T_3158 = _RAND_340[21:0];
  _RAND_341 = {1{`RANDOM}};
  _T_3097 = _RAND_341[21:0];
  _RAND_342 = {1{`RANDOM}};
  _T_3036 = _RAND_342[21:0];
  _RAND_343 = {1{`RANDOM}};
  _T_2975 = _RAND_343[21:0];
  _RAND_344 = {1{`RANDOM}};
  _T_2914 = _RAND_344[21:0];
  _RAND_345 = {1{`RANDOM}};
  _T_2853 = _RAND_345[21:0];
  _RAND_346 = {1{`RANDOM}};
  _T_2792 = _RAND_346[21:0];
  _RAND_347 = {1{`RANDOM}};
  _T_2731 = _RAND_347[21:0];
  _RAND_348 = {1{`RANDOM}};
  _T_2670 = _RAND_348[21:0];
  _RAND_349 = {1{`RANDOM}};
  _T_2609 = _RAND_349[21:0];
  _RAND_350 = {1{`RANDOM}};
  _T_2548 = _RAND_350[21:0];
  _RAND_351 = {1{`RANDOM}};
  _T_2487 = _RAND_351[21:0];
  _RAND_352 = {1{`RANDOM}};
  _T_2426 = _RAND_352[21:0];
  _RAND_353 = {1{`RANDOM}};
  _T_2365 = _RAND_353[21:0];
  _RAND_354 = {1{`RANDOM}};
  _T_2304 = _RAND_354[21:0];
  _RAND_355 = {1{`RANDOM}};
  _T_2243 = _RAND_355[21:0];
  _RAND_356 = {1{`RANDOM}};
  _T_2182 = _RAND_356[21:0];
  _RAND_357 = {1{`RANDOM}};
  _T_2121 = _RAND_357[21:0];
  _RAND_358 = {1{`RANDOM}};
  _T_2060 = _RAND_358[21:0];
  _RAND_359 = {1{`RANDOM}};
  _T_1999 = _RAND_359[21:0];
  _RAND_360 = {1{`RANDOM}};
  _T_1938 = _RAND_360[21:0];
  _RAND_361 = {1{`RANDOM}};
  _T_1877 = _RAND_361[21:0];
  _RAND_362 = {1{`RANDOM}};
  _T_1816 = _RAND_362[21:0];
  _RAND_363 = {1{`RANDOM}};
  _T_1755 = _RAND_363[21:0];
  _RAND_364 = {1{`RANDOM}};
  _T_1694 = _RAND_364[21:0];
  _RAND_365 = {1{`RANDOM}};
  _T_1633 = _RAND_365[21:0];
  _RAND_366 = {1{`RANDOM}};
  _T_1572 = _RAND_366[21:0];
  _RAND_367 = {1{`RANDOM}};
  _T_1511 = _RAND_367[21:0];
  _RAND_368 = {1{`RANDOM}};
  _T_1450 = _RAND_368[21:0];
  _RAND_369 = {1{`RANDOM}};
  _T_1389 = _RAND_369[21:0];
  _RAND_370 = {1{`RANDOM}};
  _T_1328 = _RAND_370[21:0];
  _RAND_371 = {1{`RANDOM}};
  _T_1267 = _RAND_371[21:0];
  _RAND_372 = {1{`RANDOM}};
  _T_1206 = _RAND_372[21:0];
  _RAND_373 = {1{`RANDOM}};
  _T_1145 = _RAND_373[21:0];
  _RAND_374 = {1{`RANDOM}};
  _T_1084 = _RAND_374[21:0];
  _RAND_375 = {1{`RANDOM}};
  _T_1023 = _RAND_375[21:0];
  _RAND_376 = {1{`RANDOM}};
  _T_962 = _RAND_376[21:0];
  _RAND_377 = {1{`RANDOM}};
  _T_901 = _RAND_377[21:0];
  _RAND_378 = {1{`RANDOM}};
  _T_840 = _RAND_378[21:0];
  _RAND_379 = {1{`RANDOM}};
  _T_779 = _RAND_379[21:0];
  _RAND_380 = {1{`RANDOM}};
  _T_718 = _RAND_380[21:0];
  _RAND_381 = {1{`RANDOM}};
  _T_657 = _RAND_381[21:0];
  _RAND_382 = {1{`RANDOM}};
  _T_596 = _RAND_382[21:0];
  _RAND_383 = {1{`RANDOM}};
  _T_535 = _RAND_383[21:0];
  _RAND_384 = {1{`RANDOM}};
  _T_474 = _RAND_384[21:0];
  _RAND_385 = {1{`RANDOM}};
  _T_4339 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  _T_4278 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  _T_4217 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  _T_4156 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  _T_4095 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  _T_4034 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  _T_3973 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  _T_3912 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  _T_3851 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  _T_3790 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  _T_3729 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  _T_3668 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  _T_3607 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  _T_3546 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  _T_3485 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  _T_3424 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  _T_3363 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  _T_3302 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  _T_3241 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  _T_3180 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  _T_3119 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  _T_3058 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  _T_2997 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  _T_2936 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  _T_2875 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  _T_2814 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  _T_2753 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  _T_2692 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  _T_2631 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  _T_2570 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  _T_2509 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  _T_2448 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  _T_2387 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  _T_2326 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  _T_2265 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  _T_2204 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  _T_2143 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  _T_2082 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  _T_2021 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  _T_1960 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  _T_1899 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  _T_1838 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  _T_1777 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  _T_1716 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  _T_1655 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  _T_1594 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  _T_1533 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  _T_1472 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  _T_1411 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  _T_1350 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  _T_1289 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  _T_1228 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  _T_1167 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  _T_1106 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  _T_1045 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  _T_984 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  _T_923 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  _T_862 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  _T_801 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  _T_740 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  _T_679 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  _T_618 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  _T_557 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  _T_496 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  _T_4331 = _RAND_449[21:0];
  _RAND_450 = {1{`RANDOM}};
  _T_4270 = _RAND_450[21:0];
  _RAND_451 = {1{`RANDOM}};
  _T_4209 = _RAND_451[21:0];
  _RAND_452 = {1{`RANDOM}};
  _T_4148 = _RAND_452[21:0];
  _RAND_453 = {1{`RANDOM}};
  _T_4087 = _RAND_453[21:0];
  _RAND_454 = {1{`RANDOM}};
  _T_4026 = _RAND_454[21:0];
  _RAND_455 = {1{`RANDOM}};
  _T_3965 = _RAND_455[21:0];
  _RAND_456 = {1{`RANDOM}};
  _T_3904 = _RAND_456[21:0];
  _RAND_457 = {1{`RANDOM}};
  _T_3843 = _RAND_457[21:0];
  _RAND_458 = {1{`RANDOM}};
  _T_3782 = _RAND_458[21:0];
  _RAND_459 = {1{`RANDOM}};
  _T_3721 = _RAND_459[21:0];
  _RAND_460 = {1{`RANDOM}};
  _T_3660 = _RAND_460[21:0];
  _RAND_461 = {1{`RANDOM}};
  _T_3599 = _RAND_461[21:0];
  _RAND_462 = {1{`RANDOM}};
  _T_3538 = _RAND_462[21:0];
  _RAND_463 = {1{`RANDOM}};
  _T_3477 = _RAND_463[21:0];
  _RAND_464 = {1{`RANDOM}};
  _T_3416 = _RAND_464[21:0];
  _RAND_465 = {1{`RANDOM}};
  _T_3355 = _RAND_465[21:0];
  _RAND_466 = {1{`RANDOM}};
  _T_3294 = _RAND_466[21:0];
  _RAND_467 = {1{`RANDOM}};
  _T_3233 = _RAND_467[21:0];
  _RAND_468 = {1{`RANDOM}};
  _T_3172 = _RAND_468[21:0];
  _RAND_469 = {1{`RANDOM}};
  _T_3111 = _RAND_469[21:0];
  _RAND_470 = {1{`RANDOM}};
  _T_3050 = _RAND_470[21:0];
  _RAND_471 = {1{`RANDOM}};
  _T_2989 = _RAND_471[21:0];
  _RAND_472 = {1{`RANDOM}};
  _T_2928 = _RAND_472[21:0];
  _RAND_473 = {1{`RANDOM}};
  _T_2867 = _RAND_473[21:0];
  _RAND_474 = {1{`RANDOM}};
  _T_2806 = _RAND_474[21:0];
  _RAND_475 = {1{`RANDOM}};
  _T_2745 = _RAND_475[21:0];
  _RAND_476 = {1{`RANDOM}};
  _T_2684 = _RAND_476[21:0];
  _RAND_477 = {1{`RANDOM}};
  _T_2623 = _RAND_477[21:0];
  _RAND_478 = {1{`RANDOM}};
  _T_2562 = _RAND_478[21:0];
  _RAND_479 = {1{`RANDOM}};
  _T_2501 = _RAND_479[21:0];
  _RAND_480 = {1{`RANDOM}};
  _T_2440 = _RAND_480[21:0];
  _RAND_481 = {1{`RANDOM}};
  _T_2379 = _RAND_481[21:0];
  _RAND_482 = {1{`RANDOM}};
  _T_2318 = _RAND_482[21:0];
  _RAND_483 = {1{`RANDOM}};
  _T_2257 = _RAND_483[21:0];
  _RAND_484 = {1{`RANDOM}};
  _T_2196 = _RAND_484[21:0];
  _RAND_485 = {1{`RANDOM}};
  _T_2135 = _RAND_485[21:0];
  _RAND_486 = {1{`RANDOM}};
  _T_2074 = _RAND_486[21:0];
  _RAND_487 = {1{`RANDOM}};
  _T_2013 = _RAND_487[21:0];
  _RAND_488 = {1{`RANDOM}};
  _T_1952 = _RAND_488[21:0];
  _RAND_489 = {1{`RANDOM}};
  _T_1891 = _RAND_489[21:0];
  _RAND_490 = {1{`RANDOM}};
  _T_1830 = _RAND_490[21:0];
  _RAND_491 = {1{`RANDOM}};
  _T_1769 = _RAND_491[21:0];
  _RAND_492 = {1{`RANDOM}};
  _T_1708 = _RAND_492[21:0];
  _RAND_493 = {1{`RANDOM}};
  _T_1647 = _RAND_493[21:0];
  _RAND_494 = {1{`RANDOM}};
  _T_1586 = _RAND_494[21:0];
  _RAND_495 = {1{`RANDOM}};
  _T_1525 = _RAND_495[21:0];
  _RAND_496 = {1{`RANDOM}};
  _T_1464 = _RAND_496[21:0];
  _RAND_497 = {1{`RANDOM}};
  _T_1403 = _RAND_497[21:0];
  _RAND_498 = {1{`RANDOM}};
  _T_1342 = _RAND_498[21:0];
  _RAND_499 = {1{`RANDOM}};
  _T_1281 = _RAND_499[21:0];
  _RAND_500 = {1{`RANDOM}};
  _T_1220 = _RAND_500[21:0];
  _RAND_501 = {1{`RANDOM}};
  _T_1159 = _RAND_501[21:0];
  _RAND_502 = {1{`RANDOM}};
  _T_1098 = _RAND_502[21:0];
  _RAND_503 = {1{`RANDOM}};
  _T_1037 = _RAND_503[21:0];
  _RAND_504 = {1{`RANDOM}};
  _T_976 = _RAND_504[21:0];
  _RAND_505 = {1{`RANDOM}};
  _T_915 = _RAND_505[21:0];
  _RAND_506 = {1{`RANDOM}};
  _T_854 = _RAND_506[21:0];
  _RAND_507 = {1{`RANDOM}};
  _T_793 = _RAND_507[21:0];
  _RAND_508 = {1{`RANDOM}};
  _T_732 = _RAND_508[21:0];
  _RAND_509 = {1{`RANDOM}};
  _T_671 = _RAND_509[21:0];
  _RAND_510 = {1{`RANDOM}};
  _T_610 = _RAND_510[21:0];
  _RAND_511 = {1{`RANDOM}};
  _T_549 = _RAND_511[21:0];
  _RAND_512 = {1{`RANDOM}};
  _T_488 = _RAND_512[21:0];
  _RAND_513 = {1{`RANDOM}};
  _T_501 = _RAND_513[1:0];
  _RAND_514 = {1{`RANDOM}};
  _T_440 = _RAND_514[1:0];
  _RAND_515 = {1{`RANDOM}};
  _T_562 = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  _T_623 = _RAND_516[1:0];
  _RAND_517 = {1{`RANDOM}};
  _T_684 = _RAND_517[1:0];
  _RAND_518 = {1{`RANDOM}};
  _T_745 = _RAND_518[1:0];
  _RAND_519 = {1{`RANDOM}};
  _T_806 = _RAND_519[1:0];
  _RAND_520 = {1{`RANDOM}};
  _T_867 = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  _T_928 = _RAND_521[1:0];
  _RAND_522 = {1{`RANDOM}};
  _T_989 = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  _T_1050 = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  _T_1111 = _RAND_524[1:0];
  _RAND_525 = {1{`RANDOM}};
  _T_1172 = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  _T_1233 = _RAND_526[1:0];
  _RAND_527 = {1{`RANDOM}};
  _T_1294 = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  _T_1355 = _RAND_528[1:0];
  _RAND_529 = {1{`RANDOM}};
  _T_1416 = _RAND_529[1:0];
  _RAND_530 = {1{`RANDOM}};
  _T_1477 = _RAND_530[1:0];
  _RAND_531 = {1{`RANDOM}};
  _T_1538 = _RAND_531[1:0];
  _RAND_532 = {1{`RANDOM}};
  _T_1599 = _RAND_532[1:0];
  _RAND_533 = {1{`RANDOM}};
  _T_1660 = _RAND_533[1:0];
  _RAND_534 = {1{`RANDOM}};
  _T_1721 = _RAND_534[1:0];
  _RAND_535 = {1{`RANDOM}};
  _T_1782 = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  _T_1843 = _RAND_536[1:0];
  _RAND_537 = {1{`RANDOM}};
  _T_1904 = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  _T_1965 = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  _T_2026 = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  _T_2087 = _RAND_540[1:0];
  _RAND_541 = {1{`RANDOM}};
  _T_2148 = _RAND_541[1:0];
  _RAND_542 = {1{`RANDOM}};
  _T_2209 = _RAND_542[1:0];
  _RAND_543 = {1{`RANDOM}};
  _T_2270 = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  _T_2331 = _RAND_544[1:0];
  _RAND_545 = {1{`RANDOM}};
  _T_2392 = _RAND_545[1:0];
  _RAND_546 = {1{`RANDOM}};
  _T_2453 = _RAND_546[1:0];
  _RAND_547 = {1{`RANDOM}};
  _T_2514 = _RAND_547[1:0];
  _RAND_548 = {1{`RANDOM}};
  _T_2575 = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  _T_2636 = _RAND_549[1:0];
  _RAND_550 = {1{`RANDOM}};
  _T_2697 = _RAND_550[1:0];
  _RAND_551 = {1{`RANDOM}};
  _T_2758 = _RAND_551[1:0];
  _RAND_552 = {1{`RANDOM}};
  _T_2819 = _RAND_552[1:0];
  _RAND_553 = {1{`RANDOM}};
  _T_2880 = _RAND_553[1:0];
  _RAND_554 = {1{`RANDOM}};
  _T_2941 = _RAND_554[1:0];
  _RAND_555 = {1{`RANDOM}};
  _T_3002 = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  _T_3063 = _RAND_556[1:0];
  _RAND_557 = {1{`RANDOM}};
  _T_3124 = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  _T_3185 = _RAND_558[1:0];
  _RAND_559 = {1{`RANDOM}};
  _T_3246 = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  _T_3307 = _RAND_560[1:0];
  _RAND_561 = {1{`RANDOM}};
  _T_3368 = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  _T_3429 = _RAND_562[1:0];
  _RAND_563 = {1{`RANDOM}};
  _T_3490 = _RAND_563[1:0];
  _RAND_564 = {1{`RANDOM}};
  _T_3551 = _RAND_564[1:0];
  _RAND_565 = {1{`RANDOM}};
  _T_3612 = _RAND_565[1:0];
  _RAND_566 = {1{`RANDOM}};
  _T_3673 = _RAND_566[1:0];
  _RAND_567 = {1{`RANDOM}};
  _T_3734 = _RAND_567[1:0];
  _RAND_568 = {1{`RANDOM}};
  _T_3795 = _RAND_568[1:0];
  _RAND_569 = {1{`RANDOM}};
  _T_3856 = _RAND_569[1:0];
  _RAND_570 = {1{`RANDOM}};
  _T_3917 = _RAND_570[1:0];
  _RAND_571 = {1{`RANDOM}};
  _T_3978 = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  _T_4039 = _RAND_572[1:0];
  _RAND_573 = {1{`RANDOM}};
  _T_4100 = _RAND_573[1:0];
  _RAND_574 = {1{`RANDOM}};
  _T_4161 = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  _T_4222 = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  _T_4283 = _RAND_576[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_4 <= 3'h0;
    end else if (_T_22) begin
      if (io_block) begin
        _T_4 <= 3'h4;
      end else begin
        _T_4 <= 3'h0;
      end
    end else if (_T_20) begin
      if (io_cacheOut_w_ready_i) begin
        if (io_block) begin
          _T_4 <= 3'h4;
        end else begin
          _T_4 <= 3'h0;
        end
      end else begin
        _T_4 <= 3'h3;
      end
    end else if (_T_18) begin
      if (io_block) begin
        _T_4 <= 3'h2;
      end else begin
        _T_4 <= 3'h0;
      end
    end else if (_T_16) begin
      if (io_cacheOut_r_last_i) begin
        _T_4 <= 3'h0;
      end else begin
        _T_4 <= 3'h1;
      end
    end else if (_T_14) begin
      if (io_cacheIn_valid) begin
        if (io_cacheIn_wen) begin
          _T_4 <= 3'h3;
        end else if (_T_294) begin
          _T_4 <= 3'h2;
        end else begin
          _T_4 <= 3'h1;
        end
      end else begin
        _T_4 <= 3'h0;
      end
    end else begin
      _T_4 <= 3'h0;
    end
    if (_T_448) begin
      _T_4297 <= 1'h0;
    end else begin
      _T_4297 <= _GEN_569;
    end
    if (_T_448) begin
      _T_4236 <= 1'h0;
    end else begin
      _T_4236 <= _GEN_560;
    end
    if (_T_448) begin
      _T_4175 <= 1'h0;
    end else begin
      _T_4175 <= _GEN_551;
    end
    if (_T_448) begin
      _T_4114 <= 1'h0;
    end else begin
      _T_4114 <= _GEN_542;
    end
    if (_T_448) begin
      _T_4053 <= 1'h0;
    end else begin
      _T_4053 <= _GEN_533;
    end
    if (_T_448) begin
      _T_3992 <= 1'h0;
    end else begin
      _T_3992 <= _GEN_524;
    end
    if (_T_448) begin
      _T_3931 <= 1'h0;
    end else begin
      _T_3931 <= _GEN_515;
    end
    if (_T_448) begin
      _T_3870 <= 1'h0;
    end else begin
      _T_3870 <= _GEN_506;
    end
    if (_T_448) begin
      _T_3809 <= 1'h0;
    end else begin
      _T_3809 <= _GEN_497;
    end
    if (_T_448) begin
      _T_3748 <= 1'h0;
    end else begin
      _T_3748 <= _GEN_488;
    end
    if (_T_448) begin
      _T_3687 <= 1'h0;
    end else begin
      _T_3687 <= _GEN_479;
    end
    if (_T_448) begin
      _T_3626 <= 1'h0;
    end else begin
      _T_3626 <= _GEN_470;
    end
    if (_T_448) begin
      _T_3565 <= 1'h0;
    end else begin
      _T_3565 <= _GEN_461;
    end
    if (_T_448) begin
      _T_3504 <= 1'h0;
    end else begin
      _T_3504 <= _GEN_452;
    end
    if (_T_448) begin
      _T_3443 <= 1'h0;
    end else begin
      _T_3443 <= _GEN_443;
    end
    if (_T_448) begin
      _T_3382 <= 1'h0;
    end else begin
      _T_3382 <= _GEN_434;
    end
    if (_T_448) begin
      _T_3321 <= 1'h0;
    end else begin
      _T_3321 <= _GEN_425;
    end
    if (_T_448) begin
      _T_3260 <= 1'h0;
    end else begin
      _T_3260 <= _GEN_416;
    end
    if (_T_448) begin
      _T_3199 <= 1'h0;
    end else begin
      _T_3199 <= _GEN_407;
    end
    if (_T_448) begin
      _T_3138 <= 1'h0;
    end else begin
      _T_3138 <= _GEN_398;
    end
    if (_T_448) begin
      _T_3077 <= 1'h0;
    end else begin
      _T_3077 <= _GEN_389;
    end
    if (_T_448) begin
      _T_3016 <= 1'h0;
    end else begin
      _T_3016 <= _GEN_380;
    end
    if (_T_448) begin
      _T_2955 <= 1'h0;
    end else begin
      _T_2955 <= _GEN_371;
    end
    if (_T_448) begin
      _T_2894 <= 1'h0;
    end else begin
      _T_2894 <= _GEN_362;
    end
    if (_T_448) begin
      _T_2833 <= 1'h0;
    end else begin
      _T_2833 <= _GEN_353;
    end
    if (_T_448) begin
      _T_2772 <= 1'h0;
    end else begin
      _T_2772 <= _GEN_344;
    end
    if (_T_448) begin
      _T_2711 <= 1'h0;
    end else begin
      _T_2711 <= _GEN_335;
    end
    if (_T_448) begin
      _T_2650 <= 1'h0;
    end else begin
      _T_2650 <= _GEN_326;
    end
    if (_T_448) begin
      _T_2589 <= 1'h0;
    end else begin
      _T_2589 <= _GEN_317;
    end
    if (_T_448) begin
      _T_2528 <= 1'h0;
    end else begin
      _T_2528 <= _GEN_308;
    end
    if (_T_448) begin
      _T_2467 <= 1'h0;
    end else begin
      _T_2467 <= _GEN_299;
    end
    if (_T_448) begin
      _T_2406 <= 1'h0;
    end else begin
      _T_2406 <= _GEN_290;
    end
    if (_T_448) begin
      _T_2345 <= 1'h0;
    end else begin
      _T_2345 <= _GEN_281;
    end
    if (_T_448) begin
      _T_2284 <= 1'h0;
    end else begin
      _T_2284 <= _GEN_272;
    end
    if (_T_448) begin
      _T_2223 <= 1'h0;
    end else begin
      _T_2223 <= _GEN_263;
    end
    if (_T_448) begin
      _T_2162 <= 1'h0;
    end else begin
      _T_2162 <= _GEN_254;
    end
    if (_T_448) begin
      _T_2101 <= 1'h0;
    end else begin
      _T_2101 <= _GEN_245;
    end
    if (_T_448) begin
      _T_2040 <= 1'h0;
    end else begin
      _T_2040 <= _GEN_236;
    end
    if (_T_448) begin
      _T_1979 <= 1'h0;
    end else begin
      _T_1979 <= _GEN_227;
    end
    if (_T_448) begin
      _T_1918 <= 1'h0;
    end else begin
      _T_1918 <= _GEN_218;
    end
    if (_T_448) begin
      _T_1857 <= 1'h0;
    end else begin
      _T_1857 <= _GEN_209;
    end
    if (_T_448) begin
      _T_1796 <= 1'h0;
    end else begin
      _T_1796 <= _GEN_200;
    end
    if (_T_448) begin
      _T_1735 <= 1'h0;
    end else begin
      _T_1735 <= _GEN_191;
    end
    if (_T_448) begin
      _T_1674 <= 1'h0;
    end else begin
      _T_1674 <= _GEN_182;
    end
    if (_T_448) begin
      _T_1613 <= 1'h0;
    end else begin
      _T_1613 <= _GEN_173;
    end
    if (_T_448) begin
      _T_1552 <= 1'h0;
    end else begin
      _T_1552 <= _GEN_164;
    end
    if (_T_448) begin
      _T_1491 <= 1'h0;
    end else begin
      _T_1491 <= _GEN_155;
    end
    if (_T_448) begin
      _T_1430 <= 1'h0;
    end else begin
      _T_1430 <= _GEN_146;
    end
    if (_T_448) begin
      _T_1369 <= 1'h0;
    end else begin
      _T_1369 <= _GEN_137;
    end
    if (_T_448) begin
      _T_1308 <= 1'h0;
    end else begin
      _T_1308 <= _GEN_128;
    end
    if (_T_448) begin
      _T_1247 <= 1'h0;
    end else begin
      _T_1247 <= _GEN_119;
    end
    if (_T_448) begin
      _T_1186 <= 1'h0;
    end else begin
      _T_1186 <= _GEN_110;
    end
    if (_T_448) begin
      _T_1125 <= 1'h0;
    end else begin
      _T_1125 <= _GEN_101;
    end
    if (_T_448) begin
      _T_1064 <= 1'h0;
    end else begin
      _T_1064 <= _GEN_92;
    end
    if (_T_448) begin
      _T_1003 <= 1'h0;
    end else begin
      _T_1003 <= _GEN_83;
    end
    if (_T_448) begin
      _T_942 <= 1'h0;
    end else begin
      _T_942 <= _GEN_74;
    end
    if (_T_448) begin
      _T_881 <= 1'h0;
    end else begin
      _T_881 <= _GEN_65;
    end
    if (_T_448) begin
      _T_820 <= 1'h0;
    end else begin
      _T_820 <= _GEN_56;
    end
    if (_T_448) begin
      _T_759 <= 1'h0;
    end else begin
      _T_759 <= _GEN_47;
    end
    if (_T_448) begin
      _T_698 <= 1'h0;
    end else begin
      _T_698 <= _GEN_38;
    end
    if (_T_448) begin
      _T_637 <= 1'h0;
    end else begin
      _T_637 <= _GEN_29;
    end
    if (_T_448) begin
      _T_576 <= 1'h0;
    end else begin
      _T_576 <= _GEN_20;
    end
    if (_T_448) begin
      _T_515 <= 1'h0;
    end else begin
      _T_515 <= _GEN_11;
    end
    if (_T_448) begin
      _T_454 <= 1'h0;
    end else begin
      _T_454 <= _GEN_2;
    end
    if (reset) begin
      _T_4289 <= 22'h0;
    end else if (_T_4288) begin
      _T_4289 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4228 <= 22'h0;
    end else if (_T_4227) begin
      _T_4228 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4167 <= 22'h0;
    end else if (_T_4166) begin
      _T_4167 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4106 <= 22'h0;
    end else if (_T_4105) begin
      _T_4106 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4045 <= 22'h0;
    end else if (_T_4044) begin
      _T_4045 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3984 <= 22'h0;
    end else if (_T_3983) begin
      _T_3984 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3923 <= 22'h0;
    end else if (_T_3922) begin
      _T_3923 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3862 <= 22'h0;
    end else if (_T_3861) begin
      _T_3862 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3801 <= 22'h0;
    end else if (_T_3800) begin
      _T_3801 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3740 <= 22'h0;
    end else if (_T_3739) begin
      _T_3740 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3679 <= 22'h0;
    end else if (_T_3678) begin
      _T_3679 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3618 <= 22'h0;
    end else if (_T_3617) begin
      _T_3618 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3557 <= 22'h0;
    end else if (_T_3556) begin
      _T_3557 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3496 <= 22'h0;
    end else if (_T_3495) begin
      _T_3496 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3435 <= 22'h0;
    end else if (_T_3434) begin
      _T_3435 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3374 <= 22'h0;
    end else if (_T_3373) begin
      _T_3374 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3313 <= 22'h0;
    end else if (_T_3312) begin
      _T_3313 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3252 <= 22'h0;
    end else if (_T_3251) begin
      _T_3252 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3191 <= 22'h0;
    end else if (_T_3190) begin
      _T_3191 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3130 <= 22'h0;
    end else if (_T_3129) begin
      _T_3130 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3069 <= 22'h0;
    end else if (_T_3068) begin
      _T_3069 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3008 <= 22'h0;
    end else if (_T_3007) begin
      _T_3008 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2947 <= 22'h0;
    end else if (_T_2946) begin
      _T_2947 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2886 <= 22'h0;
    end else if (_T_2885) begin
      _T_2886 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2825 <= 22'h0;
    end else if (_T_2824) begin
      _T_2825 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2764 <= 22'h0;
    end else if (_T_2763) begin
      _T_2764 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2703 <= 22'h0;
    end else if (_T_2702) begin
      _T_2703 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2642 <= 22'h0;
    end else if (_T_2641) begin
      _T_2642 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2581 <= 22'h0;
    end else if (_T_2580) begin
      _T_2581 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2520 <= 22'h0;
    end else if (_T_2519) begin
      _T_2520 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2459 <= 22'h0;
    end else if (_T_2458) begin
      _T_2459 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2398 <= 22'h0;
    end else if (_T_2397) begin
      _T_2398 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2337 <= 22'h0;
    end else if (_T_2336) begin
      _T_2337 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2276 <= 22'h0;
    end else if (_T_2275) begin
      _T_2276 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2215 <= 22'h0;
    end else if (_T_2214) begin
      _T_2215 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2154 <= 22'h0;
    end else if (_T_2153) begin
      _T_2154 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2093 <= 22'h0;
    end else if (_T_2092) begin
      _T_2093 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2032 <= 22'h0;
    end else if (_T_2031) begin
      _T_2032 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1971 <= 22'h0;
    end else if (_T_1970) begin
      _T_1971 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1910 <= 22'h0;
    end else if (_T_1909) begin
      _T_1910 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1849 <= 22'h0;
    end else if (_T_1848) begin
      _T_1849 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1788 <= 22'h0;
    end else if (_T_1787) begin
      _T_1788 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1727 <= 22'h0;
    end else if (_T_1726) begin
      _T_1727 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1666 <= 22'h0;
    end else if (_T_1665) begin
      _T_1666 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1605 <= 22'h0;
    end else if (_T_1604) begin
      _T_1605 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1544 <= 22'h0;
    end else if (_T_1543) begin
      _T_1544 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1483 <= 22'h0;
    end else if (_T_1482) begin
      _T_1483 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1422 <= 22'h0;
    end else if (_T_1421) begin
      _T_1422 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1361 <= 22'h0;
    end else if (_T_1360) begin
      _T_1361 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1300 <= 22'h0;
    end else if (_T_1299) begin
      _T_1300 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1239 <= 22'h0;
    end else if (_T_1238) begin
      _T_1239 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1178 <= 22'h0;
    end else if (_T_1177) begin
      _T_1178 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1117 <= 22'h0;
    end else if (_T_1116) begin
      _T_1117 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1056 <= 22'h0;
    end else if (_T_1055) begin
      _T_1056 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_995 <= 22'h0;
    end else if (_T_994) begin
      _T_995 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_934 <= 22'h0;
    end else if (_T_933) begin
      _T_934 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_873 <= 22'h0;
    end else if (_T_872) begin
      _T_873 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_812 <= 22'h0;
    end else if (_T_811) begin
      _T_812 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_751 <= 22'h0;
    end else if (_T_750) begin
      _T_751 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_690 <= 22'h0;
    end else if (_T_689) begin
      _T_690 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_629 <= 22'h0;
    end else if (_T_628) begin
      _T_629 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_568 <= 22'h0;
    end else if (_T_567) begin
      _T_568 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_507 <= 22'h0;
    end else if (_T_506) begin
      _T_507 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_446 <= 22'h0;
    end else if (_T_445) begin
      _T_446 <= io_cacheIn_addr[31:10];
    end
    if (_T_448) begin
      _T_4311 <= 1'h0;
    end else begin
      _T_4311 <= _GEN_571;
    end
    if (_T_448) begin
      _T_4250 <= 1'h0;
    end else begin
      _T_4250 <= _GEN_562;
    end
    if (_T_448) begin
      _T_4189 <= 1'h0;
    end else begin
      _T_4189 <= _GEN_553;
    end
    if (_T_448) begin
      _T_4128 <= 1'h0;
    end else begin
      _T_4128 <= _GEN_544;
    end
    if (_T_448) begin
      _T_4067 <= 1'h0;
    end else begin
      _T_4067 <= _GEN_535;
    end
    if (_T_448) begin
      _T_4006 <= 1'h0;
    end else begin
      _T_4006 <= _GEN_526;
    end
    if (_T_448) begin
      _T_3945 <= 1'h0;
    end else begin
      _T_3945 <= _GEN_517;
    end
    if (_T_448) begin
      _T_3884 <= 1'h0;
    end else begin
      _T_3884 <= _GEN_508;
    end
    if (_T_448) begin
      _T_3823 <= 1'h0;
    end else begin
      _T_3823 <= _GEN_499;
    end
    if (_T_448) begin
      _T_3762 <= 1'h0;
    end else begin
      _T_3762 <= _GEN_490;
    end
    if (_T_448) begin
      _T_3701 <= 1'h0;
    end else begin
      _T_3701 <= _GEN_481;
    end
    if (_T_448) begin
      _T_3640 <= 1'h0;
    end else begin
      _T_3640 <= _GEN_472;
    end
    if (_T_448) begin
      _T_3579 <= 1'h0;
    end else begin
      _T_3579 <= _GEN_463;
    end
    if (_T_448) begin
      _T_3518 <= 1'h0;
    end else begin
      _T_3518 <= _GEN_454;
    end
    if (_T_448) begin
      _T_3457 <= 1'h0;
    end else begin
      _T_3457 <= _GEN_445;
    end
    if (_T_448) begin
      _T_3396 <= 1'h0;
    end else begin
      _T_3396 <= _GEN_436;
    end
    if (_T_448) begin
      _T_3335 <= 1'h0;
    end else begin
      _T_3335 <= _GEN_427;
    end
    if (_T_448) begin
      _T_3274 <= 1'h0;
    end else begin
      _T_3274 <= _GEN_418;
    end
    if (_T_448) begin
      _T_3213 <= 1'h0;
    end else begin
      _T_3213 <= _GEN_409;
    end
    if (_T_448) begin
      _T_3152 <= 1'h0;
    end else begin
      _T_3152 <= _GEN_400;
    end
    if (_T_448) begin
      _T_3091 <= 1'h0;
    end else begin
      _T_3091 <= _GEN_391;
    end
    if (_T_448) begin
      _T_3030 <= 1'h0;
    end else begin
      _T_3030 <= _GEN_382;
    end
    if (_T_448) begin
      _T_2969 <= 1'h0;
    end else begin
      _T_2969 <= _GEN_373;
    end
    if (_T_448) begin
      _T_2908 <= 1'h0;
    end else begin
      _T_2908 <= _GEN_364;
    end
    if (_T_448) begin
      _T_2847 <= 1'h0;
    end else begin
      _T_2847 <= _GEN_355;
    end
    if (_T_448) begin
      _T_2786 <= 1'h0;
    end else begin
      _T_2786 <= _GEN_346;
    end
    if (_T_448) begin
      _T_2725 <= 1'h0;
    end else begin
      _T_2725 <= _GEN_337;
    end
    if (_T_448) begin
      _T_2664 <= 1'h0;
    end else begin
      _T_2664 <= _GEN_328;
    end
    if (_T_448) begin
      _T_2603 <= 1'h0;
    end else begin
      _T_2603 <= _GEN_319;
    end
    if (_T_448) begin
      _T_2542 <= 1'h0;
    end else begin
      _T_2542 <= _GEN_310;
    end
    if (_T_448) begin
      _T_2481 <= 1'h0;
    end else begin
      _T_2481 <= _GEN_301;
    end
    if (_T_448) begin
      _T_2420 <= 1'h0;
    end else begin
      _T_2420 <= _GEN_292;
    end
    if (_T_448) begin
      _T_2359 <= 1'h0;
    end else begin
      _T_2359 <= _GEN_283;
    end
    if (_T_448) begin
      _T_2298 <= 1'h0;
    end else begin
      _T_2298 <= _GEN_274;
    end
    if (_T_448) begin
      _T_2237 <= 1'h0;
    end else begin
      _T_2237 <= _GEN_265;
    end
    if (_T_448) begin
      _T_2176 <= 1'h0;
    end else begin
      _T_2176 <= _GEN_256;
    end
    if (_T_448) begin
      _T_2115 <= 1'h0;
    end else begin
      _T_2115 <= _GEN_247;
    end
    if (_T_448) begin
      _T_2054 <= 1'h0;
    end else begin
      _T_2054 <= _GEN_238;
    end
    if (_T_448) begin
      _T_1993 <= 1'h0;
    end else begin
      _T_1993 <= _GEN_229;
    end
    if (_T_448) begin
      _T_1932 <= 1'h0;
    end else begin
      _T_1932 <= _GEN_220;
    end
    if (_T_448) begin
      _T_1871 <= 1'h0;
    end else begin
      _T_1871 <= _GEN_211;
    end
    if (_T_448) begin
      _T_1810 <= 1'h0;
    end else begin
      _T_1810 <= _GEN_202;
    end
    if (_T_448) begin
      _T_1749 <= 1'h0;
    end else begin
      _T_1749 <= _GEN_193;
    end
    if (_T_448) begin
      _T_1688 <= 1'h0;
    end else begin
      _T_1688 <= _GEN_184;
    end
    if (_T_448) begin
      _T_1627 <= 1'h0;
    end else begin
      _T_1627 <= _GEN_175;
    end
    if (_T_448) begin
      _T_1566 <= 1'h0;
    end else begin
      _T_1566 <= _GEN_166;
    end
    if (_T_448) begin
      _T_1505 <= 1'h0;
    end else begin
      _T_1505 <= _GEN_157;
    end
    if (_T_448) begin
      _T_1444 <= 1'h0;
    end else begin
      _T_1444 <= _GEN_148;
    end
    if (_T_448) begin
      _T_1383 <= 1'h0;
    end else begin
      _T_1383 <= _GEN_139;
    end
    if (_T_448) begin
      _T_1322 <= 1'h0;
    end else begin
      _T_1322 <= _GEN_130;
    end
    if (_T_448) begin
      _T_1261 <= 1'h0;
    end else begin
      _T_1261 <= _GEN_121;
    end
    if (_T_448) begin
      _T_1200 <= 1'h0;
    end else begin
      _T_1200 <= _GEN_112;
    end
    if (_T_448) begin
      _T_1139 <= 1'h0;
    end else begin
      _T_1139 <= _GEN_103;
    end
    if (_T_448) begin
      _T_1078 <= 1'h0;
    end else begin
      _T_1078 <= _GEN_94;
    end
    if (_T_448) begin
      _T_1017 <= 1'h0;
    end else begin
      _T_1017 <= _GEN_85;
    end
    if (_T_448) begin
      _T_956 <= 1'h0;
    end else begin
      _T_956 <= _GEN_76;
    end
    if (_T_448) begin
      _T_895 <= 1'h0;
    end else begin
      _T_895 <= _GEN_67;
    end
    if (_T_448) begin
      _T_834 <= 1'h0;
    end else begin
      _T_834 <= _GEN_58;
    end
    if (_T_448) begin
      _T_773 <= 1'h0;
    end else begin
      _T_773 <= _GEN_49;
    end
    if (_T_448) begin
      _T_712 <= 1'h0;
    end else begin
      _T_712 <= _GEN_40;
    end
    if (_T_448) begin
      _T_651 <= 1'h0;
    end else begin
      _T_651 <= _GEN_31;
    end
    if (_T_448) begin
      _T_590 <= 1'h0;
    end else begin
      _T_590 <= _GEN_22;
    end
    if (_T_448) begin
      _T_529 <= 1'h0;
    end else begin
      _T_529 <= _GEN_13;
    end
    if (_T_448) begin
      _T_468 <= 1'h0;
    end else begin
      _T_468 <= _GEN_4;
    end
    if (reset) begin
      _T_4303 <= 22'h0;
    end else if (_T_4302) begin
      _T_4303 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4242 <= 22'h0;
    end else if (_T_4241) begin
      _T_4242 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4181 <= 22'h0;
    end else if (_T_4180) begin
      _T_4181 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4120 <= 22'h0;
    end else if (_T_4119) begin
      _T_4120 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4059 <= 22'h0;
    end else if (_T_4058) begin
      _T_4059 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3998 <= 22'h0;
    end else if (_T_3997) begin
      _T_3998 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3937 <= 22'h0;
    end else if (_T_3936) begin
      _T_3937 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3876 <= 22'h0;
    end else if (_T_3875) begin
      _T_3876 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3815 <= 22'h0;
    end else if (_T_3814) begin
      _T_3815 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3754 <= 22'h0;
    end else if (_T_3753) begin
      _T_3754 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3693 <= 22'h0;
    end else if (_T_3692) begin
      _T_3693 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3632 <= 22'h0;
    end else if (_T_3631) begin
      _T_3632 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3571 <= 22'h0;
    end else if (_T_3570) begin
      _T_3571 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3510 <= 22'h0;
    end else if (_T_3509) begin
      _T_3510 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3449 <= 22'h0;
    end else if (_T_3448) begin
      _T_3449 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3388 <= 22'h0;
    end else if (_T_3387) begin
      _T_3388 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3327 <= 22'h0;
    end else if (_T_3326) begin
      _T_3327 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3266 <= 22'h0;
    end else if (_T_3265) begin
      _T_3266 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3205 <= 22'h0;
    end else if (_T_3204) begin
      _T_3205 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3144 <= 22'h0;
    end else if (_T_3143) begin
      _T_3144 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3083 <= 22'h0;
    end else if (_T_3082) begin
      _T_3083 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3022 <= 22'h0;
    end else if (_T_3021) begin
      _T_3022 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2961 <= 22'h0;
    end else if (_T_2960) begin
      _T_2961 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2900 <= 22'h0;
    end else if (_T_2899) begin
      _T_2900 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2839 <= 22'h0;
    end else if (_T_2838) begin
      _T_2839 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2778 <= 22'h0;
    end else if (_T_2777) begin
      _T_2778 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2717 <= 22'h0;
    end else if (_T_2716) begin
      _T_2717 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2656 <= 22'h0;
    end else if (_T_2655) begin
      _T_2656 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2595 <= 22'h0;
    end else if (_T_2594) begin
      _T_2595 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2534 <= 22'h0;
    end else if (_T_2533) begin
      _T_2534 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2473 <= 22'h0;
    end else if (_T_2472) begin
      _T_2473 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2412 <= 22'h0;
    end else if (_T_2411) begin
      _T_2412 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2351 <= 22'h0;
    end else if (_T_2350) begin
      _T_2351 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2290 <= 22'h0;
    end else if (_T_2289) begin
      _T_2290 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2229 <= 22'h0;
    end else if (_T_2228) begin
      _T_2229 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2168 <= 22'h0;
    end else if (_T_2167) begin
      _T_2168 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2107 <= 22'h0;
    end else if (_T_2106) begin
      _T_2107 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2046 <= 22'h0;
    end else if (_T_2045) begin
      _T_2046 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1985 <= 22'h0;
    end else if (_T_1984) begin
      _T_1985 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1924 <= 22'h0;
    end else if (_T_1923) begin
      _T_1924 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1863 <= 22'h0;
    end else if (_T_1862) begin
      _T_1863 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1802 <= 22'h0;
    end else if (_T_1801) begin
      _T_1802 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1741 <= 22'h0;
    end else if (_T_1740) begin
      _T_1741 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1680 <= 22'h0;
    end else if (_T_1679) begin
      _T_1680 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1619 <= 22'h0;
    end else if (_T_1618) begin
      _T_1619 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1558 <= 22'h0;
    end else if (_T_1557) begin
      _T_1558 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1497 <= 22'h0;
    end else if (_T_1496) begin
      _T_1497 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1436 <= 22'h0;
    end else if (_T_1435) begin
      _T_1436 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1375 <= 22'h0;
    end else if (_T_1374) begin
      _T_1375 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1314 <= 22'h0;
    end else if (_T_1313) begin
      _T_1314 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1253 <= 22'h0;
    end else if (_T_1252) begin
      _T_1253 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1192 <= 22'h0;
    end else if (_T_1191) begin
      _T_1192 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1131 <= 22'h0;
    end else if (_T_1130) begin
      _T_1131 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1070 <= 22'h0;
    end else if (_T_1069) begin
      _T_1070 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1009 <= 22'h0;
    end else if (_T_1008) begin
      _T_1009 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_948 <= 22'h0;
    end else if (_T_947) begin
      _T_948 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_887 <= 22'h0;
    end else if (_T_886) begin
      _T_887 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_826 <= 22'h0;
    end else if (_T_825) begin
      _T_826 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_765 <= 22'h0;
    end else if (_T_764) begin
      _T_765 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_704 <= 22'h0;
    end else if (_T_703) begin
      _T_704 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_643 <= 22'h0;
    end else if (_T_642) begin
      _T_643 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_582 <= 22'h0;
    end else if (_T_581) begin
      _T_582 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_521 <= 22'h0;
    end else if (_T_520) begin
      _T_521 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_460 <= 22'h0;
    end else if (_T_459) begin
      _T_460 <= io_cacheIn_addr[31:10];
    end
    if (_T_448) begin
      _T_4325 <= 1'h0;
    end else begin
      _T_4325 <= _GEN_573;
    end
    if (_T_448) begin
      _T_4264 <= 1'h0;
    end else begin
      _T_4264 <= _GEN_564;
    end
    if (_T_448) begin
      _T_4203 <= 1'h0;
    end else begin
      _T_4203 <= _GEN_555;
    end
    if (_T_448) begin
      _T_4142 <= 1'h0;
    end else begin
      _T_4142 <= _GEN_546;
    end
    if (_T_448) begin
      _T_4081 <= 1'h0;
    end else begin
      _T_4081 <= _GEN_537;
    end
    if (_T_448) begin
      _T_4020 <= 1'h0;
    end else begin
      _T_4020 <= _GEN_528;
    end
    if (_T_448) begin
      _T_3959 <= 1'h0;
    end else begin
      _T_3959 <= _GEN_519;
    end
    if (_T_448) begin
      _T_3898 <= 1'h0;
    end else begin
      _T_3898 <= _GEN_510;
    end
    if (_T_448) begin
      _T_3837 <= 1'h0;
    end else begin
      _T_3837 <= _GEN_501;
    end
    if (_T_448) begin
      _T_3776 <= 1'h0;
    end else begin
      _T_3776 <= _GEN_492;
    end
    if (_T_448) begin
      _T_3715 <= 1'h0;
    end else begin
      _T_3715 <= _GEN_483;
    end
    if (_T_448) begin
      _T_3654 <= 1'h0;
    end else begin
      _T_3654 <= _GEN_474;
    end
    if (_T_448) begin
      _T_3593 <= 1'h0;
    end else begin
      _T_3593 <= _GEN_465;
    end
    if (_T_448) begin
      _T_3532 <= 1'h0;
    end else begin
      _T_3532 <= _GEN_456;
    end
    if (_T_448) begin
      _T_3471 <= 1'h0;
    end else begin
      _T_3471 <= _GEN_447;
    end
    if (_T_448) begin
      _T_3410 <= 1'h0;
    end else begin
      _T_3410 <= _GEN_438;
    end
    if (_T_448) begin
      _T_3349 <= 1'h0;
    end else begin
      _T_3349 <= _GEN_429;
    end
    if (_T_448) begin
      _T_3288 <= 1'h0;
    end else begin
      _T_3288 <= _GEN_420;
    end
    if (_T_448) begin
      _T_3227 <= 1'h0;
    end else begin
      _T_3227 <= _GEN_411;
    end
    if (_T_448) begin
      _T_3166 <= 1'h0;
    end else begin
      _T_3166 <= _GEN_402;
    end
    if (_T_448) begin
      _T_3105 <= 1'h0;
    end else begin
      _T_3105 <= _GEN_393;
    end
    if (_T_448) begin
      _T_3044 <= 1'h0;
    end else begin
      _T_3044 <= _GEN_384;
    end
    if (_T_448) begin
      _T_2983 <= 1'h0;
    end else begin
      _T_2983 <= _GEN_375;
    end
    if (_T_448) begin
      _T_2922 <= 1'h0;
    end else begin
      _T_2922 <= _GEN_366;
    end
    if (_T_448) begin
      _T_2861 <= 1'h0;
    end else begin
      _T_2861 <= _GEN_357;
    end
    if (_T_448) begin
      _T_2800 <= 1'h0;
    end else begin
      _T_2800 <= _GEN_348;
    end
    if (_T_448) begin
      _T_2739 <= 1'h0;
    end else begin
      _T_2739 <= _GEN_339;
    end
    if (_T_448) begin
      _T_2678 <= 1'h0;
    end else begin
      _T_2678 <= _GEN_330;
    end
    if (_T_448) begin
      _T_2617 <= 1'h0;
    end else begin
      _T_2617 <= _GEN_321;
    end
    if (_T_448) begin
      _T_2556 <= 1'h0;
    end else begin
      _T_2556 <= _GEN_312;
    end
    if (_T_448) begin
      _T_2495 <= 1'h0;
    end else begin
      _T_2495 <= _GEN_303;
    end
    if (_T_448) begin
      _T_2434 <= 1'h0;
    end else begin
      _T_2434 <= _GEN_294;
    end
    if (_T_448) begin
      _T_2373 <= 1'h0;
    end else begin
      _T_2373 <= _GEN_285;
    end
    if (_T_448) begin
      _T_2312 <= 1'h0;
    end else begin
      _T_2312 <= _GEN_276;
    end
    if (_T_448) begin
      _T_2251 <= 1'h0;
    end else begin
      _T_2251 <= _GEN_267;
    end
    if (_T_448) begin
      _T_2190 <= 1'h0;
    end else begin
      _T_2190 <= _GEN_258;
    end
    if (_T_448) begin
      _T_2129 <= 1'h0;
    end else begin
      _T_2129 <= _GEN_249;
    end
    if (_T_448) begin
      _T_2068 <= 1'h0;
    end else begin
      _T_2068 <= _GEN_240;
    end
    if (_T_448) begin
      _T_2007 <= 1'h0;
    end else begin
      _T_2007 <= _GEN_231;
    end
    if (_T_448) begin
      _T_1946 <= 1'h0;
    end else begin
      _T_1946 <= _GEN_222;
    end
    if (_T_448) begin
      _T_1885 <= 1'h0;
    end else begin
      _T_1885 <= _GEN_213;
    end
    if (_T_448) begin
      _T_1824 <= 1'h0;
    end else begin
      _T_1824 <= _GEN_204;
    end
    if (_T_448) begin
      _T_1763 <= 1'h0;
    end else begin
      _T_1763 <= _GEN_195;
    end
    if (_T_448) begin
      _T_1702 <= 1'h0;
    end else begin
      _T_1702 <= _GEN_186;
    end
    if (_T_448) begin
      _T_1641 <= 1'h0;
    end else begin
      _T_1641 <= _GEN_177;
    end
    if (_T_448) begin
      _T_1580 <= 1'h0;
    end else begin
      _T_1580 <= _GEN_168;
    end
    if (_T_448) begin
      _T_1519 <= 1'h0;
    end else begin
      _T_1519 <= _GEN_159;
    end
    if (_T_448) begin
      _T_1458 <= 1'h0;
    end else begin
      _T_1458 <= _GEN_150;
    end
    if (_T_448) begin
      _T_1397 <= 1'h0;
    end else begin
      _T_1397 <= _GEN_141;
    end
    if (_T_448) begin
      _T_1336 <= 1'h0;
    end else begin
      _T_1336 <= _GEN_132;
    end
    if (_T_448) begin
      _T_1275 <= 1'h0;
    end else begin
      _T_1275 <= _GEN_123;
    end
    if (_T_448) begin
      _T_1214 <= 1'h0;
    end else begin
      _T_1214 <= _GEN_114;
    end
    if (_T_448) begin
      _T_1153 <= 1'h0;
    end else begin
      _T_1153 <= _GEN_105;
    end
    if (_T_448) begin
      _T_1092 <= 1'h0;
    end else begin
      _T_1092 <= _GEN_96;
    end
    if (_T_448) begin
      _T_1031 <= 1'h0;
    end else begin
      _T_1031 <= _GEN_87;
    end
    if (_T_448) begin
      _T_970 <= 1'h0;
    end else begin
      _T_970 <= _GEN_78;
    end
    if (_T_448) begin
      _T_909 <= 1'h0;
    end else begin
      _T_909 <= _GEN_69;
    end
    if (_T_448) begin
      _T_848 <= 1'h0;
    end else begin
      _T_848 <= _GEN_60;
    end
    if (_T_448) begin
      _T_787 <= 1'h0;
    end else begin
      _T_787 <= _GEN_51;
    end
    if (_T_448) begin
      _T_726 <= 1'h0;
    end else begin
      _T_726 <= _GEN_42;
    end
    if (_T_448) begin
      _T_665 <= 1'h0;
    end else begin
      _T_665 <= _GEN_33;
    end
    if (_T_448) begin
      _T_604 <= 1'h0;
    end else begin
      _T_604 <= _GEN_24;
    end
    if (_T_448) begin
      _T_543 <= 1'h0;
    end else begin
      _T_543 <= _GEN_15;
    end
    if (_T_448) begin
      _T_482 <= 1'h0;
    end else begin
      _T_482 <= _GEN_6;
    end
    if (reset) begin
      _T_4317 <= 22'h0;
    end else if (_T_4316) begin
      _T_4317 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4256 <= 22'h0;
    end else if (_T_4255) begin
      _T_4256 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4195 <= 22'h0;
    end else if (_T_4194) begin
      _T_4195 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4134 <= 22'h0;
    end else if (_T_4133) begin
      _T_4134 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4073 <= 22'h0;
    end else if (_T_4072) begin
      _T_4073 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4012 <= 22'h0;
    end else if (_T_4011) begin
      _T_4012 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3951 <= 22'h0;
    end else if (_T_3950) begin
      _T_3951 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3890 <= 22'h0;
    end else if (_T_3889) begin
      _T_3890 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3829 <= 22'h0;
    end else if (_T_3828) begin
      _T_3829 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3768 <= 22'h0;
    end else if (_T_3767) begin
      _T_3768 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3707 <= 22'h0;
    end else if (_T_3706) begin
      _T_3707 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3646 <= 22'h0;
    end else if (_T_3645) begin
      _T_3646 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3585 <= 22'h0;
    end else if (_T_3584) begin
      _T_3585 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3524 <= 22'h0;
    end else if (_T_3523) begin
      _T_3524 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3463 <= 22'h0;
    end else if (_T_3462) begin
      _T_3463 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3402 <= 22'h0;
    end else if (_T_3401) begin
      _T_3402 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3341 <= 22'h0;
    end else if (_T_3340) begin
      _T_3341 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3280 <= 22'h0;
    end else if (_T_3279) begin
      _T_3280 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3219 <= 22'h0;
    end else if (_T_3218) begin
      _T_3219 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3158 <= 22'h0;
    end else if (_T_3157) begin
      _T_3158 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3097 <= 22'h0;
    end else if (_T_3096) begin
      _T_3097 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3036 <= 22'h0;
    end else if (_T_3035) begin
      _T_3036 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2975 <= 22'h0;
    end else if (_T_2974) begin
      _T_2975 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2914 <= 22'h0;
    end else if (_T_2913) begin
      _T_2914 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2853 <= 22'h0;
    end else if (_T_2852) begin
      _T_2853 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2792 <= 22'h0;
    end else if (_T_2791) begin
      _T_2792 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2731 <= 22'h0;
    end else if (_T_2730) begin
      _T_2731 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2670 <= 22'h0;
    end else if (_T_2669) begin
      _T_2670 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2609 <= 22'h0;
    end else if (_T_2608) begin
      _T_2609 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2548 <= 22'h0;
    end else if (_T_2547) begin
      _T_2548 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2487 <= 22'h0;
    end else if (_T_2486) begin
      _T_2487 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2426 <= 22'h0;
    end else if (_T_2425) begin
      _T_2426 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2365 <= 22'h0;
    end else if (_T_2364) begin
      _T_2365 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2304 <= 22'h0;
    end else if (_T_2303) begin
      _T_2304 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2243 <= 22'h0;
    end else if (_T_2242) begin
      _T_2243 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2182 <= 22'h0;
    end else if (_T_2181) begin
      _T_2182 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2121 <= 22'h0;
    end else if (_T_2120) begin
      _T_2121 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2060 <= 22'h0;
    end else if (_T_2059) begin
      _T_2060 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1999 <= 22'h0;
    end else if (_T_1998) begin
      _T_1999 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1938 <= 22'h0;
    end else if (_T_1937) begin
      _T_1938 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1877 <= 22'h0;
    end else if (_T_1876) begin
      _T_1877 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1816 <= 22'h0;
    end else if (_T_1815) begin
      _T_1816 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1755 <= 22'h0;
    end else if (_T_1754) begin
      _T_1755 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1694 <= 22'h0;
    end else if (_T_1693) begin
      _T_1694 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1633 <= 22'h0;
    end else if (_T_1632) begin
      _T_1633 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1572 <= 22'h0;
    end else if (_T_1571) begin
      _T_1572 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1511 <= 22'h0;
    end else if (_T_1510) begin
      _T_1511 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1450 <= 22'h0;
    end else if (_T_1449) begin
      _T_1450 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1389 <= 22'h0;
    end else if (_T_1388) begin
      _T_1389 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1328 <= 22'h0;
    end else if (_T_1327) begin
      _T_1328 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1267 <= 22'h0;
    end else if (_T_1266) begin
      _T_1267 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1206 <= 22'h0;
    end else if (_T_1205) begin
      _T_1206 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1145 <= 22'h0;
    end else if (_T_1144) begin
      _T_1145 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1084 <= 22'h0;
    end else if (_T_1083) begin
      _T_1084 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1023 <= 22'h0;
    end else if (_T_1022) begin
      _T_1023 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_962 <= 22'h0;
    end else if (_T_961) begin
      _T_962 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_901 <= 22'h0;
    end else if (_T_900) begin
      _T_901 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_840 <= 22'h0;
    end else if (_T_839) begin
      _T_840 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_779 <= 22'h0;
    end else if (_T_778) begin
      _T_779 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_718 <= 22'h0;
    end else if (_T_717) begin
      _T_718 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_657 <= 22'h0;
    end else if (_T_656) begin
      _T_657 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_596 <= 22'h0;
    end else if (_T_595) begin
      _T_596 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_535 <= 22'h0;
    end else if (_T_534) begin
      _T_535 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_474 <= 22'h0;
    end else if (_T_473) begin
      _T_474 <= io_cacheIn_addr[31:10];
    end
    if (_T_448) begin
      _T_4339 <= 1'h0;
    end else begin
      _T_4339 <= _GEN_575;
    end
    if (_T_448) begin
      _T_4278 <= 1'h0;
    end else begin
      _T_4278 <= _GEN_566;
    end
    if (_T_448) begin
      _T_4217 <= 1'h0;
    end else begin
      _T_4217 <= _GEN_557;
    end
    if (_T_448) begin
      _T_4156 <= 1'h0;
    end else begin
      _T_4156 <= _GEN_548;
    end
    if (_T_448) begin
      _T_4095 <= 1'h0;
    end else begin
      _T_4095 <= _GEN_539;
    end
    if (_T_448) begin
      _T_4034 <= 1'h0;
    end else begin
      _T_4034 <= _GEN_530;
    end
    if (_T_448) begin
      _T_3973 <= 1'h0;
    end else begin
      _T_3973 <= _GEN_521;
    end
    if (_T_448) begin
      _T_3912 <= 1'h0;
    end else begin
      _T_3912 <= _GEN_512;
    end
    if (_T_448) begin
      _T_3851 <= 1'h0;
    end else begin
      _T_3851 <= _GEN_503;
    end
    if (_T_448) begin
      _T_3790 <= 1'h0;
    end else begin
      _T_3790 <= _GEN_494;
    end
    if (_T_448) begin
      _T_3729 <= 1'h0;
    end else begin
      _T_3729 <= _GEN_485;
    end
    if (_T_448) begin
      _T_3668 <= 1'h0;
    end else begin
      _T_3668 <= _GEN_476;
    end
    if (_T_448) begin
      _T_3607 <= 1'h0;
    end else begin
      _T_3607 <= _GEN_467;
    end
    if (_T_448) begin
      _T_3546 <= 1'h0;
    end else begin
      _T_3546 <= _GEN_458;
    end
    if (_T_448) begin
      _T_3485 <= 1'h0;
    end else begin
      _T_3485 <= _GEN_449;
    end
    if (_T_448) begin
      _T_3424 <= 1'h0;
    end else begin
      _T_3424 <= _GEN_440;
    end
    if (_T_448) begin
      _T_3363 <= 1'h0;
    end else begin
      _T_3363 <= _GEN_431;
    end
    if (_T_448) begin
      _T_3302 <= 1'h0;
    end else begin
      _T_3302 <= _GEN_422;
    end
    if (_T_448) begin
      _T_3241 <= 1'h0;
    end else begin
      _T_3241 <= _GEN_413;
    end
    if (_T_448) begin
      _T_3180 <= 1'h0;
    end else begin
      _T_3180 <= _GEN_404;
    end
    if (_T_448) begin
      _T_3119 <= 1'h0;
    end else begin
      _T_3119 <= _GEN_395;
    end
    if (_T_448) begin
      _T_3058 <= 1'h0;
    end else begin
      _T_3058 <= _GEN_386;
    end
    if (_T_448) begin
      _T_2997 <= 1'h0;
    end else begin
      _T_2997 <= _GEN_377;
    end
    if (_T_448) begin
      _T_2936 <= 1'h0;
    end else begin
      _T_2936 <= _GEN_368;
    end
    if (_T_448) begin
      _T_2875 <= 1'h0;
    end else begin
      _T_2875 <= _GEN_359;
    end
    if (_T_448) begin
      _T_2814 <= 1'h0;
    end else begin
      _T_2814 <= _GEN_350;
    end
    if (_T_448) begin
      _T_2753 <= 1'h0;
    end else begin
      _T_2753 <= _GEN_341;
    end
    if (_T_448) begin
      _T_2692 <= 1'h0;
    end else begin
      _T_2692 <= _GEN_332;
    end
    if (_T_448) begin
      _T_2631 <= 1'h0;
    end else begin
      _T_2631 <= _GEN_323;
    end
    if (_T_448) begin
      _T_2570 <= 1'h0;
    end else begin
      _T_2570 <= _GEN_314;
    end
    if (_T_448) begin
      _T_2509 <= 1'h0;
    end else begin
      _T_2509 <= _GEN_305;
    end
    if (_T_448) begin
      _T_2448 <= 1'h0;
    end else begin
      _T_2448 <= _GEN_296;
    end
    if (_T_448) begin
      _T_2387 <= 1'h0;
    end else begin
      _T_2387 <= _GEN_287;
    end
    if (_T_448) begin
      _T_2326 <= 1'h0;
    end else begin
      _T_2326 <= _GEN_278;
    end
    if (_T_448) begin
      _T_2265 <= 1'h0;
    end else begin
      _T_2265 <= _GEN_269;
    end
    if (_T_448) begin
      _T_2204 <= 1'h0;
    end else begin
      _T_2204 <= _GEN_260;
    end
    if (_T_448) begin
      _T_2143 <= 1'h0;
    end else begin
      _T_2143 <= _GEN_251;
    end
    if (_T_448) begin
      _T_2082 <= 1'h0;
    end else begin
      _T_2082 <= _GEN_242;
    end
    if (_T_448) begin
      _T_2021 <= 1'h0;
    end else begin
      _T_2021 <= _GEN_233;
    end
    if (_T_448) begin
      _T_1960 <= 1'h0;
    end else begin
      _T_1960 <= _GEN_224;
    end
    if (_T_448) begin
      _T_1899 <= 1'h0;
    end else begin
      _T_1899 <= _GEN_215;
    end
    if (_T_448) begin
      _T_1838 <= 1'h0;
    end else begin
      _T_1838 <= _GEN_206;
    end
    if (_T_448) begin
      _T_1777 <= 1'h0;
    end else begin
      _T_1777 <= _GEN_197;
    end
    if (_T_448) begin
      _T_1716 <= 1'h0;
    end else begin
      _T_1716 <= _GEN_188;
    end
    if (_T_448) begin
      _T_1655 <= 1'h0;
    end else begin
      _T_1655 <= _GEN_179;
    end
    if (_T_448) begin
      _T_1594 <= 1'h0;
    end else begin
      _T_1594 <= _GEN_170;
    end
    if (_T_448) begin
      _T_1533 <= 1'h0;
    end else begin
      _T_1533 <= _GEN_161;
    end
    if (_T_448) begin
      _T_1472 <= 1'h0;
    end else begin
      _T_1472 <= _GEN_152;
    end
    if (_T_448) begin
      _T_1411 <= 1'h0;
    end else begin
      _T_1411 <= _GEN_143;
    end
    if (_T_448) begin
      _T_1350 <= 1'h0;
    end else begin
      _T_1350 <= _GEN_134;
    end
    if (_T_448) begin
      _T_1289 <= 1'h0;
    end else begin
      _T_1289 <= _GEN_125;
    end
    if (_T_448) begin
      _T_1228 <= 1'h0;
    end else begin
      _T_1228 <= _GEN_116;
    end
    if (_T_448) begin
      _T_1167 <= 1'h0;
    end else begin
      _T_1167 <= _GEN_107;
    end
    if (_T_448) begin
      _T_1106 <= 1'h0;
    end else begin
      _T_1106 <= _GEN_98;
    end
    if (_T_448) begin
      _T_1045 <= 1'h0;
    end else begin
      _T_1045 <= _GEN_89;
    end
    if (_T_448) begin
      _T_984 <= 1'h0;
    end else begin
      _T_984 <= _GEN_80;
    end
    if (_T_448) begin
      _T_923 <= 1'h0;
    end else begin
      _T_923 <= _GEN_71;
    end
    if (_T_448) begin
      _T_862 <= 1'h0;
    end else begin
      _T_862 <= _GEN_62;
    end
    if (_T_448) begin
      _T_801 <= 1'h0;
    end else begin
      _T_801 <= _GEN_53;
    end
    if (_T_448) begin
      _T_740 <= 1'h0;
    end else begin
      _T_740 <= _GEN_44;
    end
    if (_T_448) begin
      _T_679 <= 1'h0;
    end else begin
      _T_679 <= _GEN_35;
    end
    if (_T_448) begin
      _T_618 <= 1'h0;
    end else begin
      _T_618 <= _GEN_26;
    end
    if (_T_448) begin
      _T_557 <= 1'h0;
    end else begin
      _T_557 <= _GEN_17;
    end
    if (_T_448) begin
      _T_496 <= 1'h0;
    end else begin
      _T_496 <= _GEN_8;
    end
    if (reset) begin
      _T_4331 <= 22'h0;
    end else if (_T_4330) begin
      _T_4331 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4270 <= 22'h0;
    end else if (_T_4269) begin
      _T_4270 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4209 <= 22'h0;
    end else if (_T_4208) begin
      _T_4209 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4148 <= 22'h0;
    end else if (_T_4147) begin
      _T_4148 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4087 <= 22'h0;
    end else if (_T_4086) begin
      _T_4087 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_4026 <= 22'h0;
    end else if (_T_4025) begin
      _T_4026 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3965 <= 22'h0;
    end else if (_T_3964) begin
      _T_3965 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3904 <= 22'h0;
    end else if (_T_3903) begin
      _T_3904 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3843 <= 22'h0;
    end else if (_T_3842) begin
      _T_3843 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3782 <= 22'h0;
    end else if (_T_3781) begin
      _T_3782 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3721 <= 22'h0;
    end else if (_T_3720) begin
      _T_3721 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3660 <= 22'h0;
    end else if (_T_3659) begin
      _T_3660 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3599 <= 22'h0;
    end else if (_T_3598) begin
      _T_3599 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3538 <= 22'h0;
    end else if (_T_3537) begin
      _T_3538 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3477 <= 22'h0;
    end else if (_T_3476) begin
      _T_3477 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3416 <= 22'h0;
    end else if (_T_3415) begin
      _T_3416 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3355 <= 22'h0;
    end else if (_T_3354) begin
      _T_3355 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3294 <= 22'h0;
    end else if (_T_3293) begin
      _T_3294 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3233 <= 22'h0;
    end else if (_T_3232) begin
      _T_3233 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3172 <= 22'h0;
    end else if (_T_3171) begin
      _T_3172 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3111 <= 22'h0;
    end else if (_T_3110) begin
      _T_3111 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_3050 <= 22'h0;
    end else if (_T_3049) begin
      _T_3050 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2989 <= 22'h0;
    end else if (_T_2988) begin
      _T_2989 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2928 <= 22'h0;
    end else if (_T_2927) begin
      _T_2928 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2867 <= 22'h0;
    end else if (_T_2866) begin
      _T_2867 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2806 <= 22'h0;
    end else if (_T_2805) begin
      _T_2806 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2745 <= 22'h0;
    end else if (_T_2744) begin
      _T_2745 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2684 <= 22'h0;
    end else if (_T_2683) begin
      _T_2684 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2623 <= 22'h0;
    end else if (_T_2622) begin
      _T_2623 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2562 <= 22'h0;
    end else if (_T_2561) begin
      _T_2562 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2501 <= 22'h0;
    end else if (_T_2500) begin
      _T_2501 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2440 <= 22'h0;
    end else if (_T_2439) begin
      _T_2440 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2379 <= 22'h0;
    end else if (_T_2378) begin
      _T_2379 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2318 <= 22'h0;
    end else if (_T_2317) begin
      _T_2318 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2257 <= 22'h0;
    end else if (_T_2256) begin
      _T_2257 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2196 <= 22'h0;
    end else if (_T_2195) begin
      _T_2196 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2135 <= 22'h0;
    end else if (_T_2134) begin
      _T_2135 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2074 <= 22'h0;
    end else if (_T_2073) begin
      _T_2074 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_2013 <= 22'h0;
    end else if (_T_2012) begin
      _T_2013 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1952 <= 22'h0;
    end else if (_T_1951) begin
      _T_1952 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1891 <= 22'h0;
    end else if (_T_1890) begin
      _T_1891 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1830 <= 22'h0;
    end else if (_T_1829) begin
      _T_1830 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1769 <= 22'h0;
    end else if (_T_1768) begin
      _T_1769 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1708 <= 22'h0;
    end else if (_T_1707) begin
      _T_1708 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1647 <= 22'h0;
    end else if (_T_1646) begin
      _T_1647 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1586 <= 22'h0;
    end else if (_T_1585) begin
      _T_1586 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1525 <= 22'h0;
    end else if (_T_1524) begin
      _T_1525 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1464 <= 22'h0;
    end else if (_T_1463) begin
      _T_1464 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1403 <= 22'h0;
    end else if (_T_1402) begin
      _T_1403 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1342 <= 22'h0;
    end else if (_T_1341) begin
      _T_1342 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1281 <= 22'h0;
    end else if (_T_1280) begin
      _T_1281 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1220 <= 22'h0;
    end else if (_T_1219) begin
      _T_1220 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1159 <= 22'h0;
    end else if (_T_1158) begin
      _T_1159 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1098 <= 22'h0;
    end else if (_T_1097) begin
      _T_1098 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_1037 <= 22'h0;
    end else if (_T_1036) begin
      _T_1037 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_976 <= 22'h0;
    end else if (_T_975) begin
      _T_976 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_915 <= 22'h0;
    end else if (_T_914) begin
      _T_915 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_854 <= 22'h0;
    end else if (_T_853) begin
      _T_854 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_793 <= 22'h0;
    end else if (_T_792) begin
      _T_793 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_732 <= 22'h0;
    end else if (_T_731) begin
      _T_732 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_671 <= 22'h0;
    end else if (_T_670) begin
      _T_671 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_610 <= 22'h0;
    end else if (_T_609) begin
      _T_610 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_549 <= 22'h0;
    end else if (_T_548) begin
      _T_549 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_488 <= 22'h0;
    end else if (_T_487) begin
      _T_488 <= io_cacheIn_addr[31:10];
    end
    if (reset) begin
      _T_501 <= 2'h0;
    end else if (_T_500) begin
      _T_501 <= _T_498;
    end
    if (reset) begin
      _T_440 <= 2'h0;
    end else if (_T_439) begin
      _T_440 <= _T_437;
    end
    if (reset) begin
      _T_562 <= 2'h0;
    end else if (_T_561) begin
      _T_562 <= _T_559;
    end
    if (reset) begin
      _T_623 <= 2'h0;
    end else if (_T_622) begin
      _T_623 <= _T_620;
    end
    if (reset) begin
      _T_684 <= 2'h0;
    end else if (_T_683) begin
      _T_684 <= _T_681;
    end
    if (reset) begin
      _T_745 <= 2'h0;
    end else if (_T_744) begin
      _T_745 <= _T_742;
    end
    if (reset) begin
      _T_806 <= 2'h0;
    end else if (_T_805) begin
      _T_806 <= _T_803;
    end
    if (reset) begin
      _T_867 <= 2'h0;
    end else if (_T_866) begin
      _T_867 <= _T_864;
    end
    if (reset) begin
      _T_928 <= 2'h0;
    end else if (_T_927) begin
      _T_928 <= _T_925;
    end
    if (reset) begin
      _T_989 <= 2'h0;
    end else if (_T_988) begin
      _T_989 <= _T_986;
    end
    if (reset) begin
      _T_1050 <= 2'h0;
    end else if (_T_1049) begin
      _T_1050 <= _T_1047;
    end
    if (reset) begin
      _T_1111 <= 2'h0;
    end else if (_T_1110) begin
      _T_1111 <= _T_1108;
    end
    if (reset) begin
      _T_1172 <= 2'h0;
    end else if (_T_1171) begin
      _T_1172 <= _T_1169;
    end
    if (reset) begin
      _T_1233 <= 2'h0;
    end else if (_T_1232) begin
      _T_1233 <= _T_1230;
    end
    if (reset) begin
      _T_1294 <= 2'h0;
    end else if (_T_1293) begin
      _T_1294 <= _T_1291;
    end
    if (reset) begin
      _T_1355 <= 2'h0;
    end else if (_T_1354) begin
      _T_1355 <= _T_1352;
    end
    if (reset) begin
      _T_1416 <= 2'h0;
    end else if (_T_1415) begin
      _T_1416 <= _T_1413;
    end
    if (reset) begin
      _T_1477 <= 2'h0;
    end else if (_T_1476) begin
      _T_1477 <= _T_1474;
    end
    if (reset) begin
      _T_1538 <= 2'h0;
    end else if (_T_1537) begin
      _T_1538 <= _T_1535;
    end
    if (reset) begin
      _T_1599 <= 2'h0;
    end else if (_T_1598) begin
      _T_1599 <= _T_1596;
    end
    if (reset) begin
      _T_1660 <= 2'h0;
    end else if (_T_1659) begin
      _T_1660 <= _T_1657;
    end
    if (reset) begin
      _T_1721 <= 2'h0;
    end else if (_T_1720) begin
      _T_1721 <= _T_1718;
    end
    if (reset) begin
      _T_1782 <= 2'h0;
    end else if (_T_1781) begin
      _T_1782 <= _T_1779;
    end
    if (reset) begin
      _T_1843 <= 2'h0;
    end else if (_T_1842) begin
      _T_1843 <= _T_1840;
    end
    if (reset) begin
      _T_1904 <= 2'h0;
    end else if (_T_1903) begin
      _T_1904 <= _T_1901;
    end
    if (reset) begin
      _T_1965 <= 2'h0;
    end else if (_T_1964) begin
      _T_1965 <= _T_1962;
    end
    if (reset) begin
      _T_2026 <= 2'h0;
    end else if (_T_2025) begin
      _T_2026 <= _T_2023;
    end
    if (reset) begin
      _T_2087 <= 2'h0;
    end else if (_T_2086) begin
      _T_2087 <= _T_2084;
    end
    if (reset) begin
      _T_2148 <= 2'h0;
    end else if (_T_2147) begin
      _T_2148 <= _T_2145;
    end
    if (reset) begin
      _T_2209 <= 2'h0;
    end else if (_T_2208) begin
      _T_2209 <= _T_2206;
    end
    if (reset) begin
      _T_2270 <= 2'h0;
    end else if (_T_2269) begin
      _T_2270 <= _T_2267;
    end
    if (reset) begin
      _T_2331 <= 2'h0;
    end else if (_T_2330) begin
      _T_2331 <= _T_2328;
    end
    if (reset) begin
      _T_2392 <= 2'h0;
    end else if (_T_2391) begin
      _T_2392 <= _T_2389;
    end
    if (reset) begin
      _T_2453 <= 2'h0;
    end else if (_T_2452) begin
      _T_2453 <= _T_2450;
    end
    if (reset) begin
      _T_2514 <= 2'h0;
    end else if (_T_2513) begin
      _T_2514 <= _T_2511;
    end
    if (reset) begin
      _T_2575 <= 2'h0;
    end else if (_T_2574) begin
      _T_2575 <= _T_2572;
    end
    if (reset) begin
      _T_2636 <= 2'h0;
    end else if (_T_2635) begin
      _T_2636 <= _T_2633;
    end
    if (reset) begin
      _T_2697 <= 2'h0;
    end else if (_T_2696) begin
      _T_2697 <= _T_2694;
    end
    if (reset) begin
      _T_2758 <= 2'h0;
    end else if (_T_2757) begin
      _T_2758 <= _T_2755;
    end
    if (reset) begin
      _T_2819 <= 2'h0;
    end else if (_T_2818) begin
      _T_2819 <= _T_2816;
    end
    if (reset) begin
      _T_2880 <= 2'h0;
    end else if (_T_2879) begin
      _T_2880 <= _T_2877;
    end
    if (reset) begin
      _T_2941 <= 2'h0;
    end else if (_T_2940) begin
      _T_2941 <= _T_2938;
    end
    if (reset) begin
      _T_3002 <= 2'h0;
    end else if (_T_3001) begin
      _T_3002 <= _T_2999;
    end
    if (reset) begin
      _T_3063 <= 2'h0;
    end else if (_T_3062) begin
      _T_3063 <= _T_3060;
    end
    if (reset) begin
      _T_3124 <= 2'h0;
    end else if (_T_3123) begin
      _T_3124 <= _T_3121;
    end
    if (reset) begin
      _T_3185 <= 2'h0;
    end else if (_T_3184) begin
      _T_3185 <= _T_3182;
    end
    if (reset) begin
      _T_3246 <= 2'h0;
    end else if (_T_3245) begin
      _T_3246 <= _T_3243;
    end
    if (reset) begin
      _T_3307 <= 2'h0;
    end else if (_T_3306) begin
      _T_3307 <= _T_3304;
    end
    if (reset) begin
      _T_3368 <= 2'h0;
    end else if (_T_3367) begin
      _T_3368 <= _T_3365;
    end
    if (reset) begin
      _T_3429 <= 2'h0;
    end else if (_T_3428) begin
      _T_3429 <= _T_3426;
    end
    if (reset) begin
      _T_3490 <= 2'h0;
    end else if (_T_3489) begin
      _T_3490 <= _T_3487;
    end
    if (reset) begin
      _T_3551 <= 2'h0;
    end else if (_T_3550) begin
      _T_3551 <= _T_3548;
    end
    if (reset) begin
      _T_3612 <= 2'h0;
    end else if (_T_3611) begin
      _T_3612 <= _T_3609;
    end
    if (reset) begin
      _T_3673 <= 2'h0;
    end else if (_T_3672) begin
      _T_3673 <= _T_3670;
    end
    if (reset) begin
      _T_3734 <= 2'h0;
    end else if (_T_3733) begin
      _T_3734 <= _T_3731;
    end
    if (reset) begin
      _T_3795 <= 2'h0;
    end else if (_T_3794) begin
      _T_3795 <= _T_3792;
    end
    if (reset) begin
      _T_3856 <= 2'h0;
    end else if (_T_3855) begin
      _T_3856 <= _T_3853;
    end
    if (reset) begin
      _T_3917 <= 2'h0;
    end else if (_T_3916) begin
      _T_3917 <= _T_3914;
    end
    if (reset) begin
      _T_3978 <= 2'h0;
    end else if (_T_3977) begin
      _T_3978 <= _T_3975;
    end
    if (reset) begin
      _T_4039 <= 2'h0;
    end else if (_T_4038) begin
      _T_4039 <= _T_4036;
    end
    if (reset) begin
      _T_4100 <= 2'h0;
    end else if (_T_4099) begin
      _T_4100 <= _T_4097;
    end
    if (reset) begin
      _T_4161 <= 2'h0;
    end else if (_T_4160) begin
      _T_4161 <= _T_4158;
    end
    if (reset) begin
      _T_4222 <= 2'h0;
    end else if (_T_4221) begin
      _T_4222 <= _T_4219;
    end
    if (reset) begin
      _T_4283 <= 2'h0;
    end else if (_T_4282) begin
      _T_4283 <= _T_4280;
    end
  end
endmodule
module clint(
  input         clock,
  input         reset,
  input         io_clintIO_valid,
  output [63:0] io_clintIO_data_read,
  input  [63:0] io_clintIO_data_write,
  input         io_clintIO_wen,
  input  [31:0] io_clintIO_addr,
  output        intrTimeCnt_0,
  input         startTimeCnt_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtime; // @[Reg.scala 27:20]
  wire [63:0] _T_1 = mtime + 64'h1; // @[clint.scala 22:30]
  wire  _T_3 = io_clintIO_valid & io_clintIO_wen; // @[clint.scala 24:70]
  wire  _T_6 = io_clintIO_addr == 32'h2004000; // @[clint.scala 24:105]
  wire  _T_7 = _T_3 & _T_6; // @[clint.scala 24:87]
  reg [63:0] mtimecmp; // @[Reg.scala 27:20]
  wire  _T_13 = 32'h2004000 == io_clintIO_addr; // @[Mux.scala 80:60]
  wire [63:0] _T_14 = _T_13 ? mtimecmp : 64'h0; // @[Mux.scala 80:57]
  wire  _T_15 = 32'h200bff8 == io_clintIO_addr; // @[Mux.scala 80:60]
  wire  _T_17 = mtime >= mtimecmp; // @[clint.scala 38:24]
  wire  _T_18 = _T_17 & startTimeCnt_0; // @[clint.scala 38:36]
  wire  intrTimeCnt = _T_18; // @[clint.scala 37:25 clint.scala 38:15]
  assign io_clintIO_data_read = _T_15 ? mtime : _T_14; // @[clint.scala 28:24]
  assign intrTimeCnt_0 = intrTimeCnt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtime = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mtimecmp = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      mtime <= 64'h0;
    end else if (startTimeCnt_0) begin
      mtime <= _T_1;
    end
    if (reset) begin
      mtimecmp <= 64'h0;
    end else if (_T_7) begin
      mtimecmp <= io_clintIO_data_write;
    end
  end
endmodule
module mem(
  input          clock,
  input          io_memIO_cen,
  input          io_memIO_wen,
  input  [127:0] io_memIO_wdata,
  input  [5:0]   io_memIO_addr,
  input  [127:0] io_memIO_wmask,
  output [127:0] io_memIO_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [127:0] _RAND_7;
  reg [127:0] _RAND_8;
  reg [127:0] _RAND_9;
  reg [127:0] _RAND_10;
  reg [127:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [127:0] _RAND_14;
  reg [127:0] _RAND_15;
  reg [127:0] _RAND_16;
  reg [127:0] _RAND_17;
  reg [127:0] _RAND_18;
  reg [127:0] _RAND_19;
  reg [127:0] _RAND_20;
  reg [127:0] _RAND_21;
  reg [127:0] _RAND_22;
  reg [127:0] _RAND_23;
  reg [127:0] _RAND_24;
  reg [127:0] _RAND_25;
  reg [127:0] _RAND_26;
  reg [127:0] _RAND_27;
  reg [127:0] _RAND_28;
  reg [127:0] _RAND_29;
  reg [127:0] _RAND_30;
  reg [127:0] _RAND_31;
  reg [127:0] _RAND_32;
  reg [127:0] _RAND_33;
  reg [127:0] _RAND_34;
  reg [127:0] _RAND_35;
  reg [127:0] _RAND_36;
  reg [127:0] _RAND_37;
  reg [127:0] _RAND_38;
  reg [127:0] _RAND_39;
  reg [127:0] _RAND_40;
  reg [127:0] _RAND_41;
  reg [127:0] _RAND_42;
  reg [127:0] _RAND_43;
  reg [127:0] _RAND_44;
  reg [127:0] _RAND_45;
  reg [127:0] _RAND_46;
  reg [127:0] _RAND_47;
  reg [127:0] _RAND_48;
  reg [127:0] _RAND_49;
  reg [127:0] _RAND_50;
  reg [127:0] _RAND_51;
  reg [127:0] _RAND_52;
  reg [127:0] _RAND_53;
  reg [127:0] _RAND_54;
  reg [127:0] _RAND_55;
  reg [127:0] _RAND_56;
  reg [127:0] _RAND_57;
  reg [127:0] _RAND_58;
  reg [127:0] _RAND_59;
  reg [127:0] _RAND_60;
  reg [127:0] _RAND_61;
  reg [127:0] _RAND_62;
  reg [127:0] _RAND_63;
  reg [127:0] _RAND_64;
`endif // RANDOMIZE_REG_INIT
  wire  _T = ~io_memIO_cen; // @[mem.scala 15:14]
  wire [127:0] _T_2 = ~io_memIO_wmask; // @[mem.scala 16:15]
  wire  _T_3 = ~io_memIO_wen; // @[mem.scala 17:14]
  wire [127:0] _T_6 = io_memIO_wdata & _T_2; // @[mem.scala 26:47]
  reg [127:0] _T_12; // @[Reg.scala 15:16]
  wire [127:0] _T_7 = _T_12 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_8 = _T_6 | _T_7; // @[mem.scala 26:55]
  wire  _T_9 = _T & _T_3; // @[mem.scala 26:92]
  wire  _T_10 = io_memIO_addr == 6'h0; // @[mem.scala 26:116]
  wire  _T_11 = _T_9 & _T_10; // @[mem.scala 26:99]
  reg [127:0] _T_19; // @[Reg.scala 15:16]
  wire [127:0] _T_14 = _T_19 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_15 = _T_6 | _T_14; // @[mem.scala 26:55]
  wire  _T_17 = io_memIO_addr == 6'h1; // @[mem.scala 26:116]
  wire  _T_18 = _T_9 & _T_17; // @[mem.scala 26:99]
  reg [127:0] _T_26; // @[Reg.scala 15:16]
  wire [127:0] _T_21 = _T_26 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_22 = _T_6 | _T_21; // @[mem.scala 26:55]
  wire  _T_24 = io_memIO_addr == 6'h2; // @[mem.scala 26:116]
  wire  _T_25 = _T_9 & _T_24; // @[mem.scala 26:99]
  reg [127:0] _T_33; // @[Reg.scala 15:16]
  wire [127:0] _T_28 = _T_33 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_29 = _T_6 | _T_28; // @[mem.scala 26:55]
  wire  _T_31 = io_memIO_addr == 6'h3; // @[mem.scala 26:116]
  wire  _T_32 = _T_9 & _T_31; // @[mem.scala 26:99]
  reg [127:0] _T_40; // @[Reg.scala 15:16]
  wire [127:0] _T_35 = _T_40 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_36 = _T_6 | _T_35; // @[mem.scala 26:55]
  wire  _T_38 = io_memIO_addr == 6'h4; // @[mem.scala 26:116]
  wire  _T_39 = _T_9 & _T_38; // @[mem.scala 26:99]
  reg [127:0] _T_47; // @[Reg.scala 15:16]
  wire [127:0] _T_42 = _T_47 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_43 = _T_6 | _T_42; // @[mem.scala 26:55]
  wire  _T_45 = io_memIO_addr == 6'h5; // @[mem.scala 26:116]
  wire  _T_46 = _T_9 & _T_45; // @[mem.scala 26:99]
  reg [127:0] _T_54; // @[Reg.scala 15:16]
  wire [127:0] _T_49 = _T_54 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_50 = _T_6 | _T_49; // @[mem.scala 26:55]
  wire  _T_52 = io_memIO_addr == 6'h6; // @[mem.scala 26:116]
  wire  _T_53 = _T_9 & _T_52; // @[mem.scala 26:99]
  reg [127:0] _T_61; // @[Reg.scala 15:16]
  wire [127:0] _T_56 = _T_61 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_57 = _T_6 | _T_56; // @[mem.scala 26:55]
  wire  _T_59 = io_memIO_addr == 6'h7; // @[mem.scala 26:116]
  wire  _T_60 = _T_9 & _T_59; // @[mem.scala 26:99]
  reg [127:0] _T_68; // @[Reg.scala 15:16]
  wire [127:0] _T_63 = _T_68 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_64 = _T_6 | _T_63; // @[mem.scala 26:55]
  wire  _T_66 = io_memIO_addr == 6'h8; // @[mem.scala 26:116]
  wire  _T_67 = _T_9 & _T_66; // @[mem.scala 26:99]
  reg [127:0] _T_75; // @[Reg.scala 15:16]
  wire [127:0] _T_70 = _T_75 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_71 = _T_6 | _T_70; // @[mem.scala 26:55]
  wire  _T_73 = io_memIO_addr == 6'h9; // @[mem.scala 26:116]
  wire  _T_74 = _T_9 & _T_73; // @[mem.scala 26:99]
  reg [127:0] _T_82; // @[Reg.scala 15:16]
  wire [127:0] _T_77 = _T_82 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_78 = _T_6 | _T_77; // @[mem.scala 26:55]
  wire  _T_80 = io_memIO_addr == 6'ha; // @[mem.scala 26:116]
  wire  _T_81 = _T_9 & _T_80; // @[mem.scala 26:99]
  reg [127:0] _T_89; // @[Reg.scala 15:16]
  wire [127:0] _T_84 = _T_89 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_85 = _T_6 | _T_84; // @[mem.scala 26:55]
  wire  _T_87 = io_memIO_addr == 6'hb; // @[mem.scala 26:116]
  wire  _T_88 = _T_9 & _T_87; // @[mem.scala 26:99]
  reg [127:0] _T_96; // @[Reg.scala 15:16]
  wire [127:0] _T_91 = _T_96 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_92 = _T_6 | _T_91; // @[mem.scala 26:55]
  wire  _T_94 = io_memIO_addr == 6'hc; // @[mem.scala 26:116]
  wire  _T_95 = _T_9 & _T_94; // @[mem.scala 26:99]
  reg [127:0] _T_103; // @[Reg.scala 15:16]
  wire [127:0] _T_98 = _T_103 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_99 = _T_6 | _T_98; // @[mem.scala 26:55]
  wire  _T_101 = io_memIO_addr == 6'hd; // @[mem.scala 26:116]
  wire  _T_102 = _T_9 & _T_101; // @[mem.scala 26:99]
  reg [127:0] _T_110; // @[Reg.scala 15:16]
  wire [127:0] _T_105 = _T_110 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_106 = _T_6 | _T_105; // @[mem.scala 26:55]
  wire  _T_108 = io_memIO_addr == 6'he; // @[mem.scala 26:116]
  wire  _T_109 = _T_9 & _T_108; // @[mem.scala 26:99]
  reg [127:0] _T_117; // @[Reg.scala 15:16]
  wire [127:0] _T_112 = _T_117 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_113 = _T_6 | _T_112; // @[mem.scala 26:55]
  wire  _T_115 = io_memIO_addr == 6'hf; // @[mem.scala 26:116]
  wire  _T_116 = _T_9 & _T_115; // @[mem.scala 26:99]
  reg [127:0] _T_124; // @[Reg.scala 15:16]
  wire [127:0] _T_119 = _T_124 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_120 = _T_6 | _T_119; // @[mem.scala 26:55]
  wire  _T_122 = io_memIO_addr == 6'h10; // @[mem.scala 26:116]
  wire  _T_123 = _T_9 & _T_122; // @[mem.scala 26:99]
  reg [127:0] _T_131; // @[Reg.scala 15:16]
  wire [127:0] _T_126 = _T_131 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_127 = _T_6 | _T_126; // @[mem.scala 26:55]
  wire  _T_129 = io_memIO_addr == 6'h11; // @[mem.scala 26:116]
  wire  _T_130 = _T_9 & _T_129; // @[mem.scala 26:99]
  reg [127:0] _T_138; // @[Reg.scala 15:16]
  wire [127:0] _T_133 = _T_138 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_134 = _T_6 | _T_133; // @[mem.scala 26:55]
  wire  _T_136 = io_memIO_addr == 6'h12; // @[mem.scala 26:116]
  wire  _T_137 = _T_9 & _T_136; // @[mem.scala 26:99]
  reg [127:0] _T_145; // @[Reg.scala 15:16]
  wire [127:0] _T_140 = _T_145 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_141 = _T_6 | _T_140; // @[mem.scala 26:55]
  wire  _T_143 = io_memIO_addr == 6'h13; // @[mem.scala 26:116]
  wire  _T_144 = _T_9 & _T_143; // @[mem.scala 26:99]
  reg [127:0] _T_152; // @[Reg.scala 15:16]
  wire [127:0] _T_147 = _T_152 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_148 = _T_6 | _T_147; // @[mem.scala 26:55]
  wire  _T_150 = io_memIO_addr == 6'h14; // @[mem.scala 26:116]
  wire  _T_151 = _T_9 & _T_150; // @[mem.scala 26:99]
  reg [127:0] _T_159; // @[Reg.scala 15:16]
  wire [127:0] _T_154 = _T_159 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_155 = _T_6 | _T_154; // @[mem.scala 26:55]
  wire  _T_157 = io_memIO_addr == 6'h15; // @[mem.scala 26:116]
  wire  _T_158 = _T_9 & _T_157; // @[mem.scala 26:99]
  reg [127:0] _T_166; // @[Reg.scala 15:16]
  wire [127:0] _T_161 = _T_166 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_162 = _T_6 | _T_161; // @[mem.scala 26:55]
  wire  _T_164 = io_memIO_addr == 6'h16; // @[mem.scala 26:116]
  wire  _T_165 = _T_9 & _T_164; // @[mem.scala 26:99]
  reg [127:0] _T_173; // @[Reg.scala 15:16]
  wire [127:0] _T_168 = _T_173 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_169 = _T_6 | _T_168; // @[mem.scala 26:55]
  wire  _T_171 = io_memIO_addr == 6'h17; // @[mem.scala 26:116]
  wire  _T_172 = _T_9 & _T_171; // @[mem.scala 26:99]
  reg [127:0] _T_180; // @[Reg.scala 15:16]
  wire [127:0] _T_175 = _T_180 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_176 = _T_6 | _T_175; // @[mem.scala 26:55]
  wire  _T_178 = io_memIO_addr == 6'h18; // @[mem.scala 26:116]
  wire  _T_179 = _T_9 & _T_178; // @[mem.scala 26:99]
  reg [127:0] _T_187; // @[Reg.scala 15:16]
  wire [127:0] _T_182 = _T_187 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_183 = _T_6 | _T_182; // @[mem.scala 26:55]
  wire  _T_185 = io_memIO_addr == 6'h19; // @[mem.scala 26:116]
  wire  _T_186 = _T_9 & _T_185; // @[mem.scala 26:99]
  reg [127:0] _T_194; // @[Reg.scala 15:16]
  wire [127:0] _T_189 = _T_194 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_190 = _T_6 | _T_189; // @[mem.scala 26:55]
  wire  _T_192 = io_memIO_addr == 6'h1a; // @[mem.scala 26:116]
  wire  _T_193 = _T_9 & _T_192; // @[mem.scala 26:99]
  reg [127:0] _T_201; // @[Reg.scala 15:16]
  wire [127:0] _T_196 = _T_201 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_197 = _T_6 | _T_196; // @[mem.scala 26:55]
  wire  _T_199 = io_memIO_addr == 6'h1b; // @[mem.scala 26:116]
  wire  _T_200 = _T_9 & _T_199; // @[mem.scala 26:99]
  reg [127:0] _T_208; // @[Reg.scala 15:16]
  wire [127:0] _T_203 = _T_208 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_204 = _T_6 | _T_203; // @[mem.scala 26:55]
  wire  _T_206 = io_memIO_addr == 6'h1c; // @[mem.scala 26:116]
  wire  _T_207 = _T_9 & _T_206; // @[mem.scala 26:99]
  reg [127:0] _T_215; // @[Reg.scala 15:16]
  wire [127:0] _T_210 = _T_215 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_211 = _T_6 | _T_210; // @[mem.scala 26:55]
  wire  _T_213 = io_memIO_addr == 6'h1d; // @[mem.scala 26:116]
  wire  _T_214 = _T_9 & _T_213; // @[mem.scala 26:99]
  reg [127:0] _T_222; // @[Reg.scala 15:16]
  wire [127:0] _T_217 = _T_222 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_218 = _T_6 | _T_217; // @[mem.scala 26:55]
  wire  _T_220 = io_memIO_addr == 6'h1e; // @[mem.scala 26:116]
  wire  _T_221 = _T_9 & _T_220; // @[mem.scala 26:99]
  reg [127:0] _T_229; // @[Reg.scala 15:16]
  wire [127:0] _T_224 = _T_229 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_225 = _T_6 | _T_224; // @[mem.scala 26:55]
  wire  _T_227 = io_memIO_addr == 6'h1f; // @[mem.scala 26:116]
  wire  _T_228 = _T_9 & _T_227; // @[mem.scala 26:99]
  reg [127:0] _T_236; // @[Reg.scala 15:16]
  wire [127:0] _T_231 = _T_236 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_232 = _T_6 | _T_231; // @[mem.scala 26:55]
  wire  _T_234 = io_memIO_addr == 6'h20; // @[mem.scala 26:116]
  wire  _T_235 = _T_9 & _T_234; // @[mem.scala 26:99]
  reg [127:0] _T_243; // @[Reg.scala 15:16]
  wire [127:0] _T_238 = _T_243 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_239 = _T_6 | _T_238; // @[mem.scala 26:55]
  wire  _T_241 = io_memIO_addr == 6'h21; // @[mem.scala 26:116]
  wire  _T_242 = _T_9 & _T_241; // @[mem.scala 26:99]
  reg [127:0] _T_250; // @[Reg.scala 15:16]
  wire [127:0] _T_245 = _T_250 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_246 = _T_6 | _T_245; // @[mem.scala 26:55]
  wire  _T_248 = io_memIO_addr == 6'h22; // @[mem.scala 26:116]
  wire  _T_249 = _T_9 & _T_248; // @[mem.scala 26:99]
  reg [127:0] _T_257; // @[Reg.scala 15:16]
  wire [127:0] _T_252 = _T_257 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_253 = _T_6 | _T_252; // @[mem.scala 26:55]
  wire  _T_255 = io_memIO_addr == 6'h23; // @[mem.scala 26:116]
  wire  _T_256 = _T_9 & _T_255; // @[mem.scala 26:99]
  reg [127:0] _T_264; // @[Reg.scala 15:16]
  wire [127:0] _T_259 = _T_264 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_260 = _T_6 | _T_259; // @[mem.scala 26:55]
  wire  _T_262 = io_memIO_addr == 6'h24; // @[mem.scala 26:116]
  wire  _T_263 = _T_9 & _T_262; // @[mem.scala 26:99]
  reg [127:0] _T_271; // @[Reg.scala 15:16]
  wire [127:0] _T_266 = _T_271 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_267 = _T_6 | _T_266; // @[mem.scala 26:55]
  wire  _T_269 = io_memIO_addr == 6'h25; // @[mem.scala 26:116]
  wire  _T_270 = _T_9 & _T_269; // @[mem.scala 26:99]
  reg [127:0] _T_278; // @[Reg.scala 15:16]
  wire [127:0] _T_273 = _T_278 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_274 = _T_6 | _T_273; // @[mem.scala 26:55]
  wire  _T_276 = io_memIO_addr == 6'h26; // @[mem.scala 26:116]
  wire  _T_277 = _T_9 & _T_276; // @[mem.scala 26:99]
  reg [127:0] _T_285; // @[Reg.scala 15:16]
  wire [127:0] _T_280 = _T_285 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_281 = _T_6 | _T_280; // @[mem.scala 26:55]
  wire  _T_283 = io_memIO_addr == 6'h27; // @[mem.scala 26:116]
  wire  _T_284 = _T_9 & _T_283; // @[mem.scala 26:99]
  reg [127:0] _T_292; // @[Reg.scala 15:16]
  wire [127:0] _T_287 = _T_292 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_288 = _T_6 | _T_287; // @[mem.scala 26:55]
  wire  _T_290 = io_memIO_addr == 6'h28; // @[mem.scala 26:116]
  wire  _T_291 = _T_9 & _T_290; // @[mem.scala 26:99]
  reg [127:0] _T_299; // @[Reg.scala 15:16]
  wire [127:0] _T_294 = _T_299 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_295 = _T_6 | _T_294; // @[mem.scala 26:55]
  wire  _T_297 = io_memIO_addr == 6'h29; // @[mem.scala 26:116]
  wire  _T_298 = _T_9 & _T_297; // @[mem.scala 26:99]
  reg [127:0] _T_306; // @[Reg.scala 15:16]
  wire [127:0] _T_301 = _T_306 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_302 = _T_6 | _T_301; // @[mem.scala 26:55]
  wire  _T_304 = io_memIO_addr == 6'h2a; // @[mem.scala 26:116]
  wire  _T_305 = _T_9 & _T_304; // @[mem.scala 26:99]
  reg [127:0] _T_313; // @[Reg.scala 15:16]
  wire [127:0] _T_308 = _T_313 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_309 = _T_6 | _T_308; // @[mem.scala 26:55]
  wire  _T_311 = io_memIO_addr == 6'h2b; // @[mem.scala 26:116]
  wire  _T_312 = _T_9 & _T_311; // @[mem.scala 26:99]
  reg [127:0] _T_320; // @[Reg.scala 15:16]
  wire [127:0] _T_315 = _T_320 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_316 = _T_6 | _T_315; // @[mem.scala 26:55]
  wire  _T_318 = io_memIO_addr == 6'h2c; // @[mem.scala 26:116]
  wire  _T_319 = _T_9 & _T_318; // @[mem.scala 26:99]
  reg [127:0] _T_327; // @[Reg.scala 15:16]
  wire [127:0] _T_322 = _T_327 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_323 = _T_6 | _T_322; // @[mem.scala 26:55]
  wire  _T_325 = io_memIO_addr == 6'h2d; // @[mem.scala 26:116]
  wire  _T_326 = _T_9 & _T_325; // @[mem.scala 26:99]
  reg [127:0] _T_334; // @[Reg.scala 15:16]
  wire [127:0] _T_329 = _T_334 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_330 = _T_6 | _T_329; // @[mem.scala 26:55]
  wire  _T_332 = io_memIO_addr == 6'h2e; // @[mem.scala 26:116]
  wire  _T_333 = _T_9 & _T_332; // @[mem.scala 26:99]
  reg [127:0] _T_341; // @[Reg.scala 15:16]
  wire [127:0] _T_336 = _T_341 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_337 = _T_6 | _T_336; // @[mem.scala 26:55]
  wire  _T_339 = io_memIO_addr == 6'h2f; // @[mem.scala 26:116]
  wire  _T_340 = _T_9 & _T_339; // @[mem.scala 26:99]
  reg [127:0] _T_348; // @[Reg.scala 15:16]
  wire [127:0] _T_343 = _T_348 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_344 = _T_6 | _T_343; // @[mem.scala 26:55]
  wire  _T_346 = io_memIO_addr == 6'h30; // @[mem.scala 26:116]
  wire  _T_347 = _T_9 & _T_346; // @[mem.scala 26:99]
  reg [127:0] _T_355; // @[Reg.scala 15:16]
  wire [127:0] _T_350 = _T_355 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_351 = _T_6 | _T_350; // @[mem.scala 26:55]
  wire  _T_353 = io_memIO_addr == 6'h31; // @[mem.scala 26:116]
  wire  _T_354 = _T_9 & _T_353; // @[mem.scala 26:99]
  reg [127:0] _T_362; // @[Reg.scala 15:16]
  wire [127:0] _T_357 = _T_362 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_358 = _T_6 | _T_357; // @[mem.scala 26:55]
  wire  _T_360 = io_memIO_addr == 6'h32; // @[mem.scala 26:116]
  wire  _T_361 = _T_9 & _T_360; // @[mem.scala 26:99]
  reg [127:0] _T_369; // @[Reg.scala 15:16]
  wire [127:0] _T_364 = _T_369 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_365 = _T_6 | _T_364; // @[mem.scala 26:55]
  wire  _T_367 = io_memIO_addr == 6'h33; // @[mem.scala 26:116]
  wire  _T_368 = _T_9 & _T_367; // @[mem.scala 26:99]
  reg [127:0] _T_376; // @[Reg.scala 15:16]
  wire [127:0] _T_371 = _T_376 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_372 = _T_6 | _T_371; // @[mem.scala 26:55]
  wire  _T_374 = io_memIO_addr == 6'h34; // @[mem.scala 26:116]
  wire  _T_375 = _T_9 & _T_374; // @[mem.scala 26:99]
  reg [127:0] _T_383; // @[Reg.scala 15:16]
  wire [127:0] _T_378 = _T_383 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_379 = _T_6 | _T_378; // @[mem.scala 26:55]
  wire  _T_381 = io_memIO_addr == 6'h35; // @[mem.scala 26:116]
  wire  _T_382 = _T_9 & _T_381; // @[mem.scala 26:99]
  reg [127:0] _T_390; // @[Reg.scala 15:16]
  wire [127:0] _T_385 = _T_390 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_386 = _T_6 | _T_385; // @[mem.scala 26:55]
  wire  _T_388 = io_memIO_addr == 6'h36; // @[mem.scala 26:116]
  wire  _T_389 = _T_9 & _T_388; // @[mem.scala 26:99]
  reg [127:0] _T_397; // @[Reg.scala 15:16]
  wire [127:0] _T_392 = _T_397 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_393 = _T_6 | _T_392; // @[mem.scala 26:55]
  wire  _T_395 = io_memIO_addr == 6'h37; // @[mem.scala 26:116]
  wire  _T_396 = _T_9 & _T_395; // @[mem.scala 26:99]
  reg [127:0] _T_404; // @[Reg.scala 15:16]
  wire [127:0] _T_399 = _T_404 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_400 = _T_6 | _T_399; // @[mem.scala 26:55]
  wire  _T_402 = io_memIO_addr == 6'h38; // @[mem.scala 26:116]
  wire  _T_403 = _T_9 & _T_402; // @[mem.scala 26:99]
  reg [127:0] _T_411; // @[Reg.scala 15:16]
  wire [127:0] _T_406 = _T_411 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_407 = _T_6 | _T_406; // @[mem.scala 26:55]
  wire  _T_409 = io_memIO_addr == 6'h39; // @[mem.scala 26:116]
  wire  _T_410 = _T_9 & _T_409; // @[mem.scala 26:99]
  reg [127:0] _T_418; // @[Reg.scala 15:16]
  wire [127:0] _T_413 = _T_418 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_414 = _T_6 | _T_413; // @[mem.scala 26:55]
  wire  _T_416 = io_memIO_addr == 6'h3a; // @[mem.scala 26:116]
  wire  _T_417 = _T_9 & _T_416; // @[mem.scala 26:99]
  reg [127:0] _T_425; // @[Reg.scala 15:16]
  wire [127:0] _T_420 = _T_425 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_421 = _T_6 | _T_420; // @[mem.scala 26:55]
  wire  _T_423 = io_memIO_addr == 6'h3b; // @[mem.scala 26:116]
  wire  _T_424 = _T_9 & _T_423; // @[mem.scala 26:99]
  reg [127:0] _T_432; // @[Reg.scala 15:16]
  wire [127:0] _T_427 = _T_432 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_428 = _T_6 | _T_427; // @[mem.scala 26:55]
  wire  _T_430 = io_memIO_addr == 6'h3c; // @[mem.scala 26:116]
  wire  _T_431 = _T_9 & _T_430; // @[mem.scala 26:99]
  reg [127:0] _T_439; // @[Reg.scala 15:16]
  wire [127:0] _T_434 = _T_439 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_435 = _T_6 | _T_434; // @[mem.scala 26:55]
  wire  _T_437 = io_memIO_addr == 6'h3d; // @[mem.scala 26:116]
  wire  _T_438 = _T_9 & _T_437; // @[mem.scala 26:99]
  reg [127:0] _T_446; // @[Reg.scala 15:16]
  wire [127:0] _T_441 = _T_446 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_442 = _T_6 | _T_441; // @[mem.scala 26:55]
  wire  _T_444 = io_memIO_addr == 6'h3e; // @[mem.scala 26:116]
  wire  _T_445 = _T_9 & _T_444; // @[mem.scala 26:99]
  reg [127:0] _T_453; // @[Reg.scala 15:16]
  wire [127:0] _T_448 = _T_453 & io_memIO_wmask; // @[mem.scala 26:69]
  wire [127:0] _T_449 = _T_6 | _T_448; // @[mem.scala 26:55]
  wire  _T_451 = io_memIO_addr == 6'h3f; // @[mem.scala 26:116]
  wire  _T_452 = _T_9 & _T_451; // @[mem.scala 26:99]
  wire  _T_454 = 6'h1 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_456 = 6'h2 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_458 = 6'h3 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_460 = 6'h4 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_462 = 6'h5 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_464 = 6'h6 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_466 = 6'h7 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_468 = 6'h8 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_470 = 6'h9 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_472 = 6'ha == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_474 = 6'hb == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_476 = 6'hc == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_478 = 6'hd == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_480 = 6'he == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_482 = 6'hf == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_484 = 6'h10 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_486 = 6'h11 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_488 = 6'h12 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_490 = 6'h13 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_492 = 6'h14 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_494 = 6'h15 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_496 = 6'h16 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_498 = 6'h17 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_500 = 6'h18 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_502 = 6'h19 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_504 = 6'h1a == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_506 = 6'h1b == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_508 = 6'h1c == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_510 = 6'h1d == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_512 = 6'h1e == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_514 = 6'h1f == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_516 = 6'h20 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_518 = 6'h21 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_520 = 6'h22 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_522 = 6'h23 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_524 = 6'h24 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_526 = 6'h25 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_528 = 6'h26 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_530 = 6'h27 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_532 = 6'h28 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_534 = 6'h29 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_536 = 6'h2a == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_538 = 6'h2b == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_540 = 6'h2c == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_542 = 6'h2d == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_544 = 6'h2e == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_546 = 6'h2f == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_548 = 6'h30 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_550 = 6'h31 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_552 = 6'h32 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_554 = 6'h33 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_556 = 6'h34 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_558 = 6'h35 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_560 = 6'h36 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_562 = 6'h37 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_564 = 6'h38 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_566 = 6'h39 == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_568 = 6'h3a == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_570 = 6'h3b == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_572 = 6'h3c == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_574 = 6'h3d == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_576 = 6'h3e == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_578 = 6'h3f == io_memIO_addr; // @[Mux.scala 80:60]
  wire  _T_580 = _T & io_memIO_wen; // @[mem.scala 37:9]
  reg [127:0] _T_581; // @[Reg.scala 15:16]
  assign io_memIO_rdata = _T_581; // @[mem.scala 31:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  _T_12 = _RAND_0[127:0];
  _RAND_1 = {4{`RANDOM}};
  _T_19 = _RAND_1[127:0];
  _RAND_2 = {4{`RANDOM}};
  _T_26 = _RAND_2[127:0];
  _RAND_3 = {4{`RANDOM}};
  _T_33 = _RAND_3[127:0];
  _RAND_4 = {4{`RANDOM}};
  _T_40 = _RAND_4[127:0];
  _RAND_5 = {4{`RANDOM}};
  _T_47 = _RAND_5[127:0];
  _RAND_6 = {4{`RANDOM}};
  _T_54 = _RAND_6[127:0];
  _RAND_7 = {4{`RANDOM}};
  _T_61 = _RAND_7[127:0];
  _RAND_8 = {4{`RANDOM}};
  _T_68 = _RAND_8[127:0];
  _RAND_9 = {4{`RANDOM}};
  _T_75 = _RAND_9[127:0];
  _RAND_10 = {4{`RANDOM}};
  _T_82 = _RAND_10[127:0];
  _RAND_11 = {4{`RANDOM}};
  _T_89 = _RAND_11[127:0];
  _RAND_12 = {4{`RANDOM}};
  _T_96 = _RAND_12[127:0];
  _RAND_13 = {4{`RANDOM}};
  _T_103 = _RAND_13[127:0];
  _RAND_14 = {4{`RANDOM}};
  _T_110 = _RAND_14[127:0];
  _RAND_15 = {4{`RANDOM}};
  _T_117 = _RAND_15[127:0];
  _RAND_16 = {4{`RANDOM}};
  _T_124 = _RAND_16[127:0];
  _RAND_17 = {4{`RANDOM}};
  _T_131 = _RAND_17[127:0];
  _RAND_18 = {4{`RANDOM}};
  _T_138 = _RAND_18[127:0];
  _RAND_19 = {4{`RANDOM}};
  _T_145 = _RAND_19[127:0];
  _RAND_20 = {4{`RANDOM}};
  _T_152 = _RAND_20[127:0];
  _RAND_21 = {4{`RANDOM}};
  _T_159 = _RAND_21[127:0];
  _RAND_22 = {4{`RANDOM}};
  _T_166 = _RAND_22[127:0];
  _RAND_23 = {4{`RANDOM}};
  _T_173 = _RAND_23[127:0];
  _RAND_24 = {4{`RANDOM}};
  _T_180 = _RAND_24[127:0];
  _RAND_25 = {4{`RANDOM}};
  _T_187 = _RAND_25[127:0];
  _RAND_26 = {4{`RANDOM}};
  _T_194 = _RAND_26[127:0];
  _RAND_27 = {4{`RANDOM}};
  _T_201 = _RAND_27[127:0];
  _RAND_28 = {4{`RANDOM}};
  _T_208 = _RAND_28[127:0];
  _RAND_29 = {4{`RANDOM}};
  _T_215 = _RAND_29[127:0];
  _RAND_30 = {4{`RANDOM}};
  _T_222 = _RAND_30[127:0];
  _RAND_31 = {4{`RANDOM}};
  _T_229 = _RAND_31[127:0];
  _RAND_32 = {4{`RANDOM}};
  _T_236 = _RAND_32[127:0];
  _RAND_33 = {4{`RANDOM}};
  _T_243 = _RAND_33[127:0];
  _RAND_34 = {4{`RANDOM}};
  _T_250 = _RAND_34[127:0];
  _RAND_35 = {4{`RANDOM}};
  _T_257 = _RAND_35[127:0];
  _RAND_36 = {4{`RANDOM}};
  _T_264 = _RAND_36[127:0];
  _RAND_37 = {4{`RANDOM}};
  _T_271 = _RAND_37[127:0];
  _RAND_38 = {4{`RANDOM}};
  _T_278 = _RAND_38[127:0];
  _RAND_39 = {4{`RANDOM}};
  _T_285 = _RAND_39[127:0];
  _RAND_40 = {4{`RANDOM}};
  _T_292 = _RAND_40[127:0];
  _RAND_41 = {4{`RANDOM}};
  _T_299 = _RAND_41[127:0];
  _RAND_42 = {4{`RANDOM}};
  _T_306 = _RAND_42[127:0];
  _RAND_43 = {4{`RANDOM}};
  _T_313 = _RAND_43[127:0];
  _RAND_44 = {4{`RANDOM}};
  _T_320 = _RAND_44[127:0];
  _RAND_45 = {4{`RANDOM}};
  _T_327 = _RAND_45[127:0];
  _RAND_46 = {4{`RANDOM}};
  _T_334 = _RAND_46[127:0];
  _RAND_47 = {4{`RANDOM}};
  _T_341 = _RAND_47[127:0];
  _RAND_48 = {4{`RANDOM}};
  _T_348 = _RAND_48[127:0];
  _RAND_49 = {4{`RANDOM}};
  _T_355 = _RAND_49[127:0];
  _RAND_50 = {4{`RANDOM}};
  _T_362 = _RAND_50[127:0];
  _RAND_51 = {4{`RANDOM}};
  _T_369 = _RAND_51[127:0];
  _RAND_52 = {4{`RANDOM}};
  _T_376 = _RAND_52[127:0];
  _RAND_53 = {4{`RANDOM}};
  _T_383 = _RAND_53[127:0];
  _RAND_54 = {4{`RANDOM}};
  _T_390 = _RAND_54[127:0];
  _RAND_55 = {4{`RANDOM}};
  _T_397 = _RAND_55[127:0];
  _RAND_56 = {4{`RANDOM}};
  _T_404 = _RAND_56[127:0];
  _RAND_57 = {4{`RANDOM}};
  _T_411 = _RAND_57[127:0];
  _RAND_58 = {4{`RANDOM}};
  _T_418 = _RAND_58[127:0];
  _RAND_59 = {4{`RANDOM}};
  _T_425 = _RAND_59[127:0];
  _RAND_60 = {4{`RANDOM}};
  _T_432 = _RAND_60[127:0];
  _RAND_61 = {4{`RANDOM}};
  _T_439 = _RAND_61[127:0];
  _RAND_62 = {4{`RANDOM}};
  _T_446 = _RAND_62[127:0];
  _RAND_63 = {4{`RANDOM}};
  _T_453 = _RAND_63[127:0];
  _RAND_64 = {4{`RANDOM}};
  _T_581 = _RAND_64[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_11) begin
      _T_12 <= _T_8;
    end
    if (_T_18) begin
      _T_19 <= _T_15;
    end
    if (_T_25) begin
      _T_26 <= _T_22;
    end
    if (_T_32) begin
      _T_33 <= _T_29;
    end
    if (_T_39) begin
      _T_40 <= _T_36;
    end
    if (_T_46) begin
      _T_47 <= _T_43;
    end
    if (_T_53) begin
      _T_54 <= _T_50;
    end
    if (_T_60) begin
      _T_61 <= _T_57;
    end
    if (_T_67) begin
      _T_68 <= _T_64;
    end
    if (_T_74) begin
      _T_75 <= _T_71;
    end
    if (_T_81) begin
      _T_82 <= _T_78;
    end
    if (_T_88) begin
      _T_89 <= _T_85;
    end
    if (_T_95) begin
      _T_96 <= _T_92;
    end
    if (_T_102) begin
      _T_103 <= _T_99;
    end
    if (_T_109) begin
      _T_110 <= _T_106;
    end
    if (_T_116) begin
      _T_117 <= _T_113;
    end
    if (_T_123) begin
      _T_124 <= _T_120;
    end
    if (_T_130) begin
      _T_131 <= _T_127;
    end
    if (_T_137) begin
      _T_138 <= _T_134;
    end
    if (_T_144) begin
      _T_145 <= _T_141;
    end
    if (_T_151) begin
      _T_152 <= _T_148;
    end
    if (_T_158) begin
      _T_159 <= _T_155;
    end
    if (_T_165) begin
      _T_166 <= _T_162;
    end
    if (_T_172) begin
      _T_173 <= _T_169;
    end
    if (_T_179) begin
      _T_180 <= _T_176;
    end
    if (_T_186) begin
      _T_187 <= _T_183;
    end
    if (_T_193) begin
      _T_194 <= _T_190;
    end
    if (_T_200) begin
      _T_201 <= _T_197;
    end
    if (_T_207) begin
      _T_208 <= _T_204;
    end
    if (_T_214) begin
      _T_215 <= _T_211;
    end
    if (_T_221) begin
      _T_222 <= _T_218;
    end
    if (_T_228) begin
      _T_229 <= _T_225;
    end
    if (_T_235) begin
      _T_236 <= _T_232;
    end
    if (_T_242) begin
      _T_243 <= _T_239;
    end
    if (_T_249) begin
      _T_250 <= _T_246;
    end
    if (_T_256) begin
      _T_257 <= _T_253;
    end
    if (_T_263) begin
      _T_264 <= _T_260;
    end
    if (_T_270) begin
      _T_271 <= _T_267;
    end
    if (_T_277) begin
      _T_278 <= _T_274;
    end
    if (_T_284) begin
      _T_285 <= _T_281;
    end
    if (_T_291) begin
      _T_292 <= _T_288;
    end
    if (_T_298) begin
      _T_299 <= _T_295;
    end
    if (_T_305) begin
      _T_306 <= _T_302;
    end
    if (_T_312) begin
      _T_313 <= _T_309;
    end
    if (_T_319) begin
      _T_320 <= _T_316;
    end
    if (_T_326) begin
      _T_327 <= _T_323;
    end
    if (_T_333) begin
      _T_334 <= _T_330;
    end
    if (_T_340) begin
      _T_341 <= _T_337;
    end
    if (_T_347) begin
      _T_348 <= _T_344;
    end
    if (_T_354) begin
      _T_355 <= _T_351;
    end
    if (_T_361) begin
      _T_362 <= _T_358;
    end
    if (_T_368) begin
      _T_369 <= _T_365;
    end
    if (_T_375) begin
      _T_376 <= _T_372;
    end
    if (_T_382) begin
      _T_383 <= _T_379;
    end
    if (_T_389) begin
      _T_390 <= _T_386;
    end
    if (_T_396) begin
      _T_397 <= _T_393;
    end
    if (_T_403) begin
      _T_404 <= _T_400;
    end
    if (_T_410) begin
      _T_411 <= _T_407;
    end
    if (_T_417) begin
      _T_418 <= _T_414;
    end
    if (_T_424) begin
      _T_425 <= _T_421;
    end
    if (_T_431) begin
      _T_432 <= _T_428;
    end
    if (_T_438) begin
      _T_439 <= _T_435;
    end
    if (_T_445) begin
      _T_446 <= _T_442;
    end
    if (_T_452) begin
      _T_453 <= _T_449;
    end
    if (_T_580) begin
      if (_T_578) begin
        _T_581 <= _T_453;
      end else if (_T_576) begin
        _T_581 <= _T_446;
      end else if (_T_574) begin
        _T_581 <= _T_439;
      end else if (_T_572) begin
        _T_581 <= _T_432;
      end else if (_T_570) begin
        _T_581 <= _T_425;
      end else if (_T_568) begin
        _T_581 <= _T_418;
      end else if (_T_566) begin
        _T_581 <= _T_411;
      end else if (_T_564) begin
        _T_581 <= _T_404;
      end else if (_T_562) begin
        _T_581 <= _T_397;
      end else if (_T_560) begin
        _T_581 <= _T_390;
      end else if (_T_558) begin
        _T_581 <= _T_383;
      end else if (_T_556) begin
        _T_581 <= _T_376;
      end else if (_T_554) begin
        _T_581 <= _T_369;
      end else if (_T_552) begin
        _T_581 <= _T_362;
      end else if (_T_550) begin
        _T_581 <= _T_355;
      end else if (_T_548) begin
        _T_581 <= _T_348;
      end else if (_T_546) begin
        _T_581 <= _T_341;
      end else if (_T_544) begin
        _T_581 <= _T_334;
      end else if (_T_542) begin
        _T_581 <= _T_327;
      end else if (_T_540) begin
        _T_581 <= _T_320;
      end else if (_T_538) begin
        _T_581 <= _T_313;
      end else if (_T_536) begin
        _T_581 <= _T_306;
      end else if (_T_534) begin
        _T_581 <= _T_299;
      end else if (_T_532) begin
        _T_581 <= _T_292;
      end else if (_T_530) begin
        _T_581 <= _T_285;
      end else if (_T_528) begin
        _T_581 <= _T_278;
      end else if (_T_526) begin
        _T_581 <= _T_271;
      end else if (_T_524) begin
        _T_581 <= _T_264;
      end else if (_T_522) begin
        _T_581 <= _T_257;
      end else if (_T_520) begin
        _T_581 <= _T_250;
      end else if (_T_518) begin
        _T_581 <= _T_243;
      end else if (_T_516) begin
        _T_581 <= _T_236;
      end else if (_T_514) begin
        _T_581 <= _T_229;
      end else if (_T_512) begin
        _T_581 <= _T_222;
      end else if (_T_510) begin
        _T_581 <= _T_215;
      end else if (_T_508) begin
        _T_581 <= _T_208;
      end else if (_T_506) begin
        _T_581 <= _T_201;
      end else if (_T_504) begin
        _T_581 <= _T_194;
      end else if (_T_502) begin
        _T_581 <= _T_187;
      end else if (_T_500) begin
        _T_581 <= _T_180;
      end else if (_T_498) begin
        _T_581 <= _T_173;
      end else if (_T_496) begin
        _T_581 <= _T_166;
      end else if (_T_494) begin
        _T_581 <= _T_159;
      end else if (_T_492) begin
        _T_581 <= _T_152;
      end else if (_T_490) begin
        _T_581 <= _T_145;
      end else if (_T_488) begin
        _T_581 <= _T_138;
      end else if (_T_486) begin
        _T_581 <= _T_131;
      end else if (_T_484) begin
        _T_581 <= _T_124;
      end else if (_T_482) begin
        _T_581 <= _T_117;
      end else if (_T_480) begin
        _T_581 <= _T_110;
      end else if (_T_478) begin
        _T_581 <= _T_103;
      end else if (_T_476) begin
        _T_581 <= _T_96;
      end else if (_T_474) begin
        _T_581 <= _T_89;
      end else if (_T_472) begin
        _T_581 <= _T_82;
      end else if (_T_470) begin
        _T_581 <= _T_75;
      end else if (_T_468) begin
        _T_581 <= _T_68;
      end else if (_T_466) begin
        _T_581 <= _T_61;
      end else if (_T_464) begin
        _T_581 <= _T_54;
      end else if (_T_462) begin
        _T_581 <= _T_47;
      end else if (_T_460) begin
        _T_581 <= _T_40;
      end else if (_T_458) begin
        _T_581 <= _T_33;
      end else if (_T_456) begin
        _T_581 <= _T_26;
      end else if (_T_454) begin
        _T_581 <= _T_19;
      end else begin
        _T_581 <= _T_12;
      end
    end
  end
endmodule
module TopOK(
  input         clock,
  input         reset,
  input         io_dmaster_awready,
  output        io_dmaster_awvalid,
  output [3:0]  io_dmaster_awid,
  output [31:0] io_dmaster_awaddr,
  output [7:0]  io_dmaster_awlen,
  output [2:0]  io_dmaster_awsize,
  output [1:0]  io_dmaster_awburst,
  input         io_dmaster_wready,
  output        io_dmaster_wvalid,
  output [63:0] io_dmaster_wdata,
  output [7:0]  io_dmaster_wstrb,
  output        io_dmaster_wlast,
  output        io_dmaster_bready,
  input         io_dmaster_bvalid,
  input  [3:0]  io_dmaster_bid,
  input  [1:0]  io_dmaster_bresp,
  input         io_dmaster_arready,
  output        io_dmaster_arvalid,
  output [3:0]  io_dmaster_arid,
  output [31:0] io_dmaster_araddr,
  output [7:0]  io_dmaster_arlen,
  output [2:0]  io_dmaster_arsize,
  output [1:0]  io_dmaster_arburst,
  output        io_dmaster_rready,
  input         io_dmaster_rvalid,
  input  [3:0]  io_dmaster_rid,
  input  [1:0]  io_dmaster_rresp,
  input  [63:0] io_dmaster_rdata,
  input         io_dmaster_rlast,
  output [32:0] io_outputs_0,
  output [32:0] io_outputs_1,
  output [32:0] io_outputs_2,
  output [32:0] io_outputs_3,
  output [32:0] io_outputs_4,
  output [32:0] io_outputs_5,
  output [32:0] io_outputs_6,
  output [32:0] io_outputs_7,
  output [32:0] io_outputs_8,
  output [32:0] io_outputs_9,
  output [32:0] io_outputs_10,
  output [32:0] io_outputs_11,
  output [32:0] io_outputs_12,
  output [32:0] io_outputs_13,
  output [32:0] io_outputs_14,
  output [32:0] io_outputs_15,
  output        io_mmio_valid,
  input         io_mmio_ready,
  input  [63:0] io_mmio_data_read,
  output [63:0] io_mmio_data_write,
  output        io_mmio_wen,
  output [31:0] io_mmio_addr,
  output [1:0]  io_mmio_rsize,
  output [7:0]  io_mmio_mask
);
  wire  dmaIns_clock; // @[Top.scala 33:22]
  wire  dmaIns_reset; // @[Top.scala 33:22]
  wire  dmaIns_io_dataIn_awready; // @[Top.scala 33:22]
  wire  dmaIns_io_dataIn_awvalid; // @[Top.scala 33:22]
  wire [31:0] dmaIns_io_dataIn_awaddr; // @[Top.scala 33:22]
  wire [7:0] dmaIns_io_dataIn_awlen; // @[Top.scala 33:22]
  wire  dmaIns_io_dataIn_wready; // @[Top.scala 33:22]
  wire  dmaIns_io_dataIn_wvalid; // @[Top.scala 33:22]
  wire [63:0] dmaIns_io_dataIn_wdata; // @[Top.scala 33:22]
  wire  dmaIns_io_dataIn_wlast; // @[Top.scala 33:22]
  wire  dmaIns_io_dataIn_bready; // @[Top.scala 33:22]
  wire  dmaIns_io_dataIn_bvalid; // @[Top.scala 33:22]
  wire  dmaIns_io_dataIn_arready; // @[Top.scala 33:22]
  wire  dmaIns_io_dataIn_arvalid; // @[Top.scala 33:22]
  wire [31:0] dmaIns_io_dataIn_araddr; // @[Top.scala 33:22]
  wire [7:0] dmaIns_io_dataIn_arlen; // @[Top.scala 33:22]
  wire  dmaIns_io_dataIn_rready; // @[Top.scala 33:22]
  wire  dmaIns_io_dataIn_rvalid; // @[Top.scala 33:22]
  wire [63:0] dmaIns_io_dataIn_rdata; // @[Top.scala 33:22]
  wire  dmaIns_io_dataIn_rlast; // @[Top.scala 33:22]
  wire  dmaIns_io_dataOutMMIO_valid; // @[Top.scala 33:22]
  wire  dmaIns_io_dataOutMMIO_ready; // @[Top.scala 33:22]
  wire [63:0] dmaIns_io_dataOutMMIO_data_read; // @[Top.scala 33:22]
  wire [63:0] dmaIns_io_dataOutMMIO_data_write; // @[Top.scala 33:22]
  wire  dmaIns_io_dataOutMMIO_wen; // @[Top.scala 33:22]
  wire [31:0] dmaIns_io_dataOutMMIO_addr; // @[Top.scala 33:22]
  wire  dmaIns_dmaEn_0; // @[Top.scala 33:22]
  wire  dmaIns_dmaEnWR_0; // @[Top.scala 33:22]
  wire  dmaIns_block3_0; // @[Top.scala 33:22]
  wire [191:0] dmaIns_dmaCtrl_0; // @[Top.scala 33:22]
  wire  dmaIns_block2_0; // @[Top.scala 33:22]
  wire  dmaIns_blockDMA_0; // @[Top.scala 33:22]
  wire  dmaIns_DMABuzy_0; // @[Top.scala 33:22]
  wire  cgraIns_clock; // @[Top.scala 34:23]
  wire  cgraIns_reset; // @[Top.scala 34:23]
  wire  cgraIns_io_CGRAIO_valid; // @[Top.scala 34:23]
  wire  cgraIns_io_CGRAIO_ready; // @[Top.scala 34:23]
  wire [63:0] cgraIns_io_CGRAIO_data_read; // @[Top.scala 34:23]
  wire [63:0] cgraIns_io_CGRAIO_data_write; // @[Top.scala 34:23]
  wire  cgraIns_io_CGRAIO_wen; // @[Top.scala 34:23]
  wire [31:0] cgraIns_io_CGRAIO_addr; // @[Top.scala 34:23]
  wire [32:0] cgraIns_io_outputs_0; // @[Top.scala 34:23]
  wire [32:0] cgraIns_io_outputs_1; // @[Top.scala 34:23]
  wire [32:0] cgraIns_io_outputs_2; // @[Top.scala 34:23]
  wire [32:0] cgraIns_io_outputs_3; // @[Top.scala 34:23]
  wire [32:0] cgraIns_io_outputs_4; // @[Top.scala 34:23]
  wire [32:0] cgraIns_io_outputs_5; // @[Top.scala 34:23]
  wire [32:0] cgraIns_io_outputs_6; // @[Top.scala 34:23]
  wire [32:0] cgraIns_io_outputs_7; // @[Top.scala 34:23]
  wire [32:0] cgraIns_io_outputs_8; // @[Top.scala 34:23]
  wire [32:0] cgraIns_io_outputs_9; // @[Top.scala 34:23]
  wire [32:0] cgraIns_io_outputs_10; // @[Top.scala 34:23]
  wire [32:0] cgraIns_io_outputs_11; // @[Top.scala 34:23]
  wire [32:0] cgraIns_io_outputs_12; // @[Top.scala 34:23]
  wire [32:0] cgraIns_io_outputs_13; // @[Top.scala 34:23]
  wire [32:0] cgraIns_io_outputs_14; // @[Top.scala 34:23]
  wire [32:0] cgraIns_io_outputs_15; // @[Top.scala 34:23]
  wire  cgraIns__T_100_0; // @[Top.scala 34:23]
  wire [191:0] cgraIns_dmaCtrl; // @[Top.scala 34:23]
  wire  riscvIns_clock; // @[Top.scala 35:24]
  wire  riscvIns_reset; // @[Top.scala 35:24]
  wire  riscvIns_io_instIO_valid; // @[Top.scala 35:24]
  wire  riscvIns_io_instIO_ready; // @[Top.scala 35:24]
  wire [63:0] riscvIns_io_instIO_data_read; // @[Top.scala 35:24]
  wire [31:0] riscvIns_io_instIO_addr; // @[Top.scala 35:24]
  wire  riscvIns_io_dataIO_valid; // @[Top.scala 35:24]
  wire  riscvIns_io_dataIO_ready; // @[Top.scala 35:24]
  wire [63:0] riscvIns_io_dataIO_data_read; // @[Top.scala 35:24]
  wire [63:0] riscvIns_io_dataIO_data_write; // @[Top.scala 35:24]
  wire  riscvIns_io_dataIO_wen; // @[Top.scala 35:24]
  wire [31:0] riscvIns_io_dataIO_addr; // @[Top.scala 35:24]
  wire [1:0] riscvIns_io_dataIO_rsize; // @[Top.scala 35:24]
  wire [7:0] riscvIns_io_dataIO_mask; // @[Top.scala 35:24]
  wire  riscvIns__T_99_0; // @[Top.scala 35:24]
  wire  riscvIns_intrTimeCnt_0; // @[Top.scala 35:24]
  wire  riscvIns__T_100_0; // @[Top.scala 35:24]
  wire  riscvIns_startTimeCnt; // @[Top.scala 35:24]
  wire  riscvIns_block3_0; // @[Top.scala 35:24]
  wire [191:0] riscvIns_dmaCtrl; // @[Top.scala 35:24]
  wire  riscvIns_block2_0; // @[Top.scala 35:24]
  wire  riscvIns_blockDMA_0; // @[Top.scala 35:24]
  wire  riscvIns_fencei_0; // @[Top.scala 35:24]
  wire  iCache_clock; // @[Top.scala 36:22]
  wire  iCache_reset; // @[Top.scala 36:22]
  wire  iCache_io_cacheOut_ar_valid_o; // @[Top.scala 36:22]
  wire [31:0] iCache_io_cacheOut_ar_addr_o; // @[Top.scala 36:22]
  wire [7:0] iCache_io_cacheOut_ar_len_o; // @[Top.scala 36:22]
  wire  iCache_io_cacheOut_r_valid_i; // @[Top.scala 36:22]
  wire [63:0] iCache_io_cacheOut_r_data_i; // @[Top.scala 36:22]
  wire  iCache_io_cacheOut_r_last_i; // @[Top.scala 36:22]
  wire [31:0] iCache_io_cacheOut_w_addr_o; // @[Top.scala 36:22]
  wire  iCache_io_cacheIn_valid; // @[Top.scala 36:22]
  wire  iCache_io_cacheIn_ready; // @[Top.scala 36:22]
  wire [63:0] iCache_io_cacheIn_data_read; // @[Top.scala 36:22]
  wire [31:0] iCache_io_cacheIn_addr; // @[Top.scala 36:22]
  wire  iCache_io_SRAMIO_0_cen; // @[Top.scala 36:22]
  wire  iCache_io_SRAMIO_0_wen; // @[Top.scala 36:22]
  wire [127:0] iCache_io_SRAMIO_0_wdata; // @[Top.scala 36:22]
  wire [5:0] iCache_io_SRAMIO_0_addr; // @[Top.scala 36:22]
  wire [127:0] iCache_io_SRAMIO_0_wmask; // @[Top.scala 36:22]
  wire [127:0] iCache_io_SRAMIO_0_rdata; // @[Top.scala 36:22]
  wire  iCache_io_SRAMIO_1_cen; // @[Top.scala 36:22]
  wire  iCache_io_SRAMIO_1_wen; // @[Top.scala 36:22]
  wire [127:0] iCache_io_SRAMIO_1_wdata; // @[Top.scala 36:22]
  wire [5:0] iCache_io_SRAMIO_1_addr; // @[Top.scala 36:22]
  wire [127:0] iCache_io_SRAMIO_1_wmask; // @[Top.scala 36:22]
  wire [127:0] iCache_io_SRAMIO_1_rdata; // @[Top.scala 36:22]
  wire  iCache_io_SRAMIO_2_cen; // @[Top.scala 36:22]
  wire  iCache_io_SRAMIO_2_wen; // @[Top.scala 36:22]
  wire [127:0] iCache_io_SRAMIO_2_wdata; // @[Top.scala 36:22]
  wire [5:0] iCache_io_SRAMIO_2_addr; // @[Top.scala 36:22]
  wire [127:0] iCache_io_SRAMIO_2_wmask; // @[Top.scala 36:22]
  wire [127:0] iCache_io_SRAMIO_2_rdata; // @[Top.scala 36:22]
  wire  iCache_io_SRAMIO_3_cen; // @[Top.scala 36:22]
  wire  iCache_io_SRAMIO_3_wen; // @[Top.scala 36:22]
  wire [127:0] iCache_io_SRAMIO_3_wdata; // @[Top.scala 36:22]
  wire [5:0] iCache_io_SRAMIO_3_addr; // @[Top.scala 36:22]
  wire [127:0] iCache_io_SRAMIO_3_wmask; // @[Top.scala 36:22]
  wire [127:0] iCache_io_SRAMIO_3_rdata; // @[Top.scala 36:22]
  wire  iCache_io_block; // @[Top.scala 36:22]
  wire  iCache_updataICache; // @[Top.scala 36:22]
  wire  axiIIO_clock; // @[Top.scala 38:22]
  wire  axiIIO_reset; // @[Top.scala 38:22]
  wire  axiIIO_io_axiIO_awready; // @[Top.scala 38:22]
  wire  axiIIO_io_axiIO_awvalid; // @[Top.scala 38:22]
  wire [31:0] axiIIO_io_axiIO_awaddr; // @[Top.scala 38:22]
  wire [2:0] axiIIO_io_axiIO_awsize; // @[Top.scala 38:22]
  wire  axiIIO_io_axiIO_wready; // @[Top.scala 38:22]
  wire  axiIIO_io_axiIO_wvalid; // @[Top.scala 38:22]
  wire [63:0] axiIIO_io_axiIO_wdata; // @[Top.scala 38:22]
  wire [7:0] axiIIO_io_axiIO_wstrb; // @[Top.scala 38:22]
  wire  axiIIO_io_axiIO_wlast; // @[Top.scala 38:22]
  wire  axiIIO_io_axiIO_bready; // @[Top.scala 38:22]
  wire  axiIIO_io_axiIO_bvalid; // @[Top.scala 38:22]
  wire  axiIIO_io_axiIO_arready; // @[Top.scala 38:22]
  wire  axiIIO_io_axiIO_arvalid; // @[Top.scala 38:22]
  wire [31:0] axiIIO_io_axiIO_araddr; // @[Top.scala 38:22]
  wire [7:0] axiIIO_io_axiIO_arlen; // @[Top.scala 38:22]
  wire [2:0] axiIIO_io_axiIO_arsize; // @[Top.scala 38:22]
  wire [1:0] axiIIO_io_axiIO_arburst; // @[Top.scala 38:22]
  wire  axiIIO_io_axiIO_rready; // @[Top.scala 38:22]
  wire  axiIIO_io_axiIO_rvalid; // @[Top.scala 38:22]
  wire [63:0] axiIIO_io_axiIO_rdata; // @[Top.scala 38:22]
  wire  axiIIO_io_axiIO_rlast; // @[Top.scala 38:22]
  wire  axiIIO_io_cache_ar_valid_o; // @[Top.scala 38:22]
  wire [31:0] axiIIO_io_cache_ar_addr_o; // @[Top.scala 38:22]
  wire [7:0] axiIIO_io_cache_ar_len_o; // @[Top.scala 38:22]
  wire  axiIIO_io_cache_r_valid_i; // @[Top.scala 38:22]
  wire [63:0] axiIIO_io_cache_r_data_i; // @[Top.scala 38:22]
  wire  axiIIO_io_cache_r_last_i; // @[Top.scala 38:22]
  wire  axiIIO_io_cache_w_valid_o; // @[Top.scala 38:22]
  wire  axiIIO_io_cache_w_ready_i; // @[Top.scala 38:22]
  wire [63:0] axiIIO_io_cache_w_data_o; // @[Top.scala 38:22]
  wire [31:0] axiIIO_io_cache_w_addr_o; // @[Top.scala 38:22]
  wire [7:0] axiIIO_io_cache_w_mask_o; // @[Top.scala 38:22]
  wire [1:0] axiIIO_io_cache_wsize; // @[Top.scala 38:22]
  wire  dArbIns_io_arbIn_valid; // @[Top.scala 41:23]
  wire  dArbIns_io_arbIn_ready; // @[Top.scala 41:23]
  wire [63:0] dArbIns_io_arbIn_data_read; // @[Top.scala 41:23]
  wire [63:0] dArbIns_io_arbIn_data_write; // @[Top.scala 41:23]
  wire  dArbIns_io_arbIn_wen; // @[Top.scala 41:23]
  wire [31:0] dArbIns_io_arbIn_addr; // @[Top.scala 41:23]
  wire [1:0] dArbIns_io_arbIn_rsize; // @[Top.scala 41:23]
  wire [7:0] dArbIns_io_arbIn_mask; // @[Top.scala 41:23]
  wire  dArbIns_io_arbMMIO_valid; // @[Top.scala 41:23]
  wire  dArbIns_io_arbMMIO_ready; // @[Top.scala 41:23]
  wire [63:0] dArbIns_io_arbMMIO_data_read; // @[Top.scala 41:23]
  wire [63:0] dArbIns_io_arbMMIO_data_write; // @[Top.scala 41:23]
  wire  dArbIns_io_arbMMIO_wen; // @[Top.scala 41:23]
  wire [31:0] dArbIns_io_arbMMIO_addr; // @[Top.scala 41:23]
  wire [1:0] dArbIns_io_arbMMIO_rsize; // @[Top.scala 41:23]
  wire [7:0] dArbIns_io_arbMMIO_mask; // @[Top.scala 41:23]
  wire  dArbIns_io_arbClint_valid; // @[Top.scala 41:23]
  wire [63:0] dArbIns_io_arbClint_data_read; // @[Top.scala 41:23]
  wire [63:0] dArbIns_io_arbClint_data_write; // @[Top.scala 41:23]
  wire  dArbIns_io_arbClint_wen; // @[Top.scala 41:23]
  wire [31:0] dArbIns_io_arbClint_addr; // @[Top.scala 41:23]
  wire  dArbIns_io_arbDCache_valid; // @[Top.scala 41:23]
  wire  dArbIns_io_arbDCache_ready; // @[Top.scala 41:23]
  wire [63:0] dArbIns_io_arbDCache_data_read; // @[Top.scala 41:23]
  wire [63:0] dArbIns_io_arbDCache_data_write; // @[Top.scala 41:23]
  wire  dArbIns_io_arbDCache_wen; // @[Top.scala 41:23]
  wire [31:0] dArbIns_io_arbDCache_addr; // @[Top.scala 41:23]
  wire [1:0] dArbIns_io_arbDCache_rsize; // @[Top.scala 41:23]
  wire [7:0] dArbIns_io_arbDCache_mask; // @[Top.scala 41:23]
  wire  dArbIns_io_arbCgra_valid; // @[Top.scala 41:23]
  wire  dArbIns_io_arbCgra_ready; // @[Top.scala 41:23]
  wire [63:0] dArbIns_io_arbCgra_data_read; // @[Top.scala 41:23]
  wire [63:0] dArbIns_io_arbCgra_data_write; // @[Top.scala 41:23]
  wire  dArbIns_io_arbCgra_wen; // @[Top.scala 41:23]
  wire [31:0] dArbIns_io_arbCgra_addr; // @[Top.scala 41:23]
  wire  mmioDCache_io_mmioIn_valid; // @[Top.scala 42:26]
  wire  mmioDCache_io_mmioIn_ready; // @[Top.scala 42:26]
  wire [63:0] mmioDCache_io_mmioIn_data_read; // @[Top.scala 42:26]
  wire [63:0] mmioDCache_io_mmioIn_data_write; // @[Top.scala 42:26]
  wire  mmioDCache_io_mmioIn_wen; // @[Top.scala 42:26]
  wire [31:0] mmioDCache_io_mmioIn_addr; // @[Top.scala 42:26]
  wire  mmioDCache_io_mmioOut_valid; // @[Top.scala 42:26]
  wire  mmioDCache_io_mmioOut_ready; // @[Top.scala 42:26]
  wire [63:0] mmioDCache_io_mmioOut_data_read; // @[Top.scala 42:26]
  wire [63:0] mmioDCache_io_mmioOut_data_write; // @[Top.scala 42:26]
  wire  mmioDCache_io_mmioOut_wen; // @[Top.scala 42:26]
  wire [31:0] mmioDCache_io_mmioOut_addr; // @[Top.scala 42:26]
  wire  dCache_clock; // @[Top.scala 43:22]
  wire  dCache_reset; // @[Top.scala 43:22]
  wire  dCache_io_cacheOut_ar_valid_o; // @[Top.scala 43:22]
  wire [31:0] dCache_io_cacheOut_ar_addr_o; // @[Top.scala 43:22]
  wire [7:0] dCache_io_cacheOut_ar_len_o; // @[Top.scala 43:22]
  wire  dCache_io_cacheOut_r_valid_i; // @[Top.scala 43:22]
  wire [63:0] dCache_io_cacheOut_r_data_i; // @[Top.scala 43:22]
  wire  dCache_io_cacheOut_r_last_i; // @[Top.scala 43:22]
  wire  dCache_io_cacheOut_w_valid_o; // @[Top.scala 43:22]
  wire  dCache_io_cacheOut_w_ready_i; // @[Top.scala 43:22]
  wire [63:0] dCache_io_cacheOut_w_data_o; // @[Top.scala 43:22]
  wire [31:0] dCache_io_cacheOut_w_addr_o; // @[Top.scala 43:22]
  wire [7:0] dCache_io_cacheOut_w_mask_o; // @[Top.scala 43:22]
  wire [1:0] dCache_io_cacheOut_wsize; // @[Top.scala 43:22]
  wire  dCache_io_cacheIn_valid; // @[Top.scala 43:22]
  wire  dCache_io_cacheIn_ready; // @[Top.scala 43:22]
  wire [63:0] dCache_io_cacheIn_data_read; // @[Top.scala 43:22]
  wire [63:0] dCache_io_cacheIn_data_write; // @[Top.scala 43:22]
  wire  dCache_io_cacheIn_wen; // @[Top.scala 43:22]
  wire [31:0] dCache_io_cacheIn_addr; // @[Top.scala 43:22]
  wire [1:0] dCache_io_cacheIn_rsize; // @[Top.scala 43:22]
  wire [7:0] dCache_io_cacheIn_mask; // @[Top.scala 43:22]
  wire  dCache_io_SRAMIO_0_cen; // @[Top.scala 43:22]
  wire  dCache_io_SRAMIO_0_wen; // @[Top.scala 43:22]
  wire [127:0] dCache_io_SRAMIO_0_wdata; // @[Top.scala 43:22]
  wire [5:0] dCache_io_SRAMIO_0_addr; // @[Top.scala 43:22]
  wire [127:0] dCache_io_SRAMIO_0_wmask; // @[Top.scala 43:22]
  wire [127:0] dCache_io_SRAMIO_0_rdata; // @[Top.scala 43:22]
  wire  dCache_io_SRAMIO_1_cen; // @[Top.scala 43:22]
  wire  dCache_io_SRAMIO_1_wen; // @[Top.scala 43:22]
  wire [127:0] dCache_io_SRAMIO_1_wdata; // @[Top.scala 43:22]
  wire [5:0] dCache_io_SRAMIO_1_addr; // @[Top.scala 43:22]
  wire [127:0] dCache_io_SRAMIO_1_wmask; // @[Top.scala 43:22]
  wire [127:0] dCache_io_SRAMIO_1_rdata; // @[Top.scala 43:22]
  wire  dCache_io_SRAMIO_2_cen; // @[Top.scala 43:22]
  wire  dCache_io_SRAMIO_2_wen; // @[Top.scala 43:22]
  wire [127:0] dCache_io_SRAMIO_2_wdata; // @[Top.scala 43:22]
  wire [5:0] dCache_io_SRAMIO_2_addr; // @[Top.scala 43:22]
  wire [127:0] dCache_io_SRAMIO_2_wmask; // @[Top.scala 43:22]
  wire [127:0] dCache_io_SRAMIO_2_rdata; // @[Top.scala 43:22]
  wire  dCache_io_SRAMIO_3_cen; // @[Top.scala 43:22]
  wire  dCache_io_SRAMIO_3_wen; // @[Top.scala 43:22]
  wire [127:0] dCache_io_SRAMIO_3_wdata; // @[Top.scala 43:22]
  wire [5:0] dCache_io_SRAMIO_3_addr; // @[Top.scala 43:22]
  wire [127:0] dCache_io_SRAMIO_3_wmask; // @[Top.scala 43:22]
  wire [127:0] dCache_io_SRAMIO_3_rdata; // @[Top.scala 43:22]
  wire  dCache_io_block; // @[Top.scala 43:22]
  wire  dCache_updataICache; // @[Top.scala 43:22]
  wire  clintIns_clock; // @[Top.scala 44:25]
  wire  clintIns_reset; // @[Top.scala 44:25]
  wire  clintIns_io_clintIO_valid; // @[Top.scala 44:25]
  wire [63:0] clintIns_io_clintIO_data_read; // @[Top.scala 44:25]
  wire [63:0] clintIns_io_clintIO_data_write; // @[Top.scala 44:25]
  wire  clintIns_io_clintIO_wen; // @[Top.scala 44:25]
  wire [31:0] clintIns_io_clintIO_addr; // @[Top.scala 44:25]
  wire  clintIns_intrTimeCnt_0; // @[Top.scala 44:25]
  wire  clintIns_startTimeCnt_0; // @[Top.scala 44:25]
  wire  axiDIO_clock; // @[Top.scala 53:22]
  wire  axiDIO_reset; // @[Top.scala 53:22]
  wire  axiDIO_io_axiIO_awready; // @[Top.scala 53:22]
  wire  axiDIO_io_axiIO_awvalid; // @[Top.scala 53:22]
  wire [31:0] axiDIO_io_axiIO_awaddr; // @[Top.scala 53:22]
  wire [2:0] axiDIO_io_axiIO_awsize; // @[Top.scala 53:22]
  wire  axiDIO_io_axiIO_wready; // @[Top.scala 53:22]
  wire  axiDIO_io_axiIO_wvalid; // @[Top.scala 53:22]
  wire [63:0] axiDIO_io_axiIO_wdata; // @[Top.scala 53:22]
  wire [7:0] axiDIO_io_axiIO_wstrb; // @[Top.scala 53:22]
  wire  axiDIO_io_axiIO_wlast; // @[Top.scala 53:22]
  wire  axiDIO_io_axiIO_bready; // @[Top.scala 53:22]
  wire  axiDIO_io_axiIO_bvalid; // @[Top.scala 53:22]
  wire  axiDIO_io_axiIO_arready; // @[Top.scala 53:22]
  wire  axiDIO_io_axiIO_arvalid; // @[Top.scala 53:22]
  wire [31:0] axiDIO_io_axiIO_araddr; // @[Top.scala 53:22]
  wire [7:0] axiDIO_io_axiIO_arlen; // @[Top.scala 53:22]
  wire [2:0] axiDIO_io_axiIO_arsize; // @[Top.scala 53:22]
  wire [1:0] axiDIO_io_axiIO_arburst; // @[Top.scala 53:22]
  wire  axiDIO_io_axiIO_rready; // @[Top.scala 53:22]
  wire  axiDIO_io_axiIO_rvalid; // @[Top.scala 53:22]
  wire [63:0] axiDIO_io_axiIO_rdata; // @[Top.scala 53:22]
  wire  axiDIO_io_axiIO_rlast; // @[Top.scala 53:22]
  wire  axiDIO_io_cache_ar_valid_o; // @[Top.scala 53:22]
  wire [31:0] axiDIO_io_cache_ar_addr_o; // @[Top.scala 53:22]
  wire [7:0] axiDIO_io_cache_ar_len_o; // @[Top.scala 53:22]
  wire  axiDIO_io_cache_r_valid_i; // @[Top.scala 53:22]
  wire [63:0] axiDIO_io_cache_r_data_i; // @[Top.scala 53:22]
  wire  axiDIO_io_cache_r_last_i; // @[Top.scala 53:22]
  wire  axiDIO_io_cache_w_valid_o; // @[Top.scala 53:22]
  wire  axiDIO_io_cache_w_ready_i; // @[Top.scala 53:22]
  wire [63:0] axiDIO_io_cache_w_data_o; // @[Top.scala 53:22]
  wire [31:0] axiDIO_io_cache_w_addr_o; // @[Top.scala 53:22]
  wire [7:0] axiDIO_io_cache_w_mask_o; // @[Top.scala 53:22]
  wire [1:0] axiDIO_io_cache_wsize; // @[Top.scala 53:22]
  wire  mem_clock; // @[Top.scala 60:24]
  wire  mem_io_memIO_cen; // @[Top.scala 60:24]
  wire  mem_io_memIO_wen; // @[Top.scala 60:24]
  wire [127:0] mem_io_memIO_wdata; // @[Top.scala 60:24]
  wire [5:0] mem_io_memIO_addr; // @[Top.scala 60:24]
  wire [127:0] mem_io_memIO_wmask; // @[Top.scala 60:24]
  wire [127:0] mem_io_memIO_rdata; // @[Top.scala 60:24]
  wire  mem_1_clock; // @[Top.scala 61:24]
  wire  mem_1_io_memIO_cen; // @[Top.scala 61:24]
  wire  mem_1_io_memIO_wen; // @[Top.scala 61:24]
  wire [127:0] mem_1_io_memIO_wdata; // @[Top.scala 61:24]
  wire [5:0] mem_1_io_memIO_addr; // @[Top.scala 61:24]
  wire [127:0] mem_1_io_memIO_wmask; // @[Top.scala 61:24]
  wire [127:0] mem_1_io_memIO_rdata; // @[Top.scala 61:24]
  wire  mem_2_clock; // @[Top.scala 60:24]
  wire  mem_2_io_memIO_cen; // @[Top.scala 60:24]
  wire  mem_2_io_memIO_wen; // @[Top.scala 60:24]
  wire [127:0] mem_2_io_memIO_wdata; // @[Top.scala 60:24]
  wire [5:0] mem_2_io_memIO_addr; // @[Top.scala 60:24]
  wire [127:0] mem_2_io_memIO_wmask; // @[Top.scala 60:24]
  wire [127:0] mem_2_io_memIO_rdata; // @[Top.scala 60:24]
  wire  mem_3_clock; // @[Top.scala 61:24]
  wire  mem_3_io_memIO_cen; // @[Top.scala 61:24]
  wire  mem_3_io_memIO_wen; // @[Top.scala 61:24]
  wire [127:0] mem_3_io_memIO_wdata; // @[Top.scala 61:24]
  wire [5:0] mem_3_io_memIO_addr; // @[Top.scala 61:24]
  wire [127:0] mem_3_io_memIO_wmask; // @[Top.scala 61:24]
  wire [127:0] mem_3_io_memIO_rdata; // @[Top.scala 61:24]
  wire  mem_4_clock; // @[Top.scala 60:24]
  wire  mem_4_io_memIO_cen; // @[Top.scala 60:24]
  wire  mem_4_io_memIO_wen; // @[Top.scala 60:24]
  wire [127:0] mem_4_io_memIO_wdata; // @[Top.scala 60:24]
  wire [5:0] mem_4_io_memIO_addr; // @[Top.scala 60:24]
  wire [127:0] mem_4_io_memIO_wmask; // @[Top.scala 60:24]
  wire [127:0] mem_4_io_memIO_rdata; // @[Top.scala 60:24]
  wire  mem_5_clock; // @[Top.scala 61:24]
  wire  mem_5_io_memIO_cen; // @[Top.scala 61:24]
  wire  mem_5_io_memIO_wen; // @[Top.scala 61:24]
  wire [127:0] mem_5_io_memIO_wdata; // @[Top.scala 61:24]
  wire [5:0] mem_5_io_memIO_addr; // @[Top.scala 61:24]
  wire [127:0] mem_5_io_memIO_wmask; // @[Top.scala 61:24]
  wire [127:0] mem_5_io_memIO_rdata; // @[Top.scala 61:24]
  wire  mem_6_clock; // @[Top.scala 60:24]
  wire  mem_6_io_memIO_cen; // @[Top.scala 60:24]
  wire  mem_6_io_memIO_wen; // @[Top.scala 60:24]
  wire [127:0] mem_6_io_memIO_wdata; // @[Top.scala 60:24]
  wire [5:0] mem_6_io_memIO_addr; // @[Top.scala 60:24]
  wire [127:0] mem_6_io_memIO_wmask; // @[Top.scala 60:24]
  wire [127:0] mem_6_io_memIO_rdata; // @[Top.scala 60:24]
  wire  mem_7_clock; // @[Top.scala 61:24]
  wire  mem_7_io_memIO_cen; // @[Top.scala 61:24]
  wire  mem_7_io_memIO_wen; // @[Top.scala 61:24]
  wire [127:0] mem_7_io_memIO_wdata; // @[Top.scala 61:24]
  wire [5:0] mem_7_io_memIO_addr; // @[Top.scala 61:24]
  wire [127:0] mem_7_io_memIO_wmask; // @[Top.scala 61:24]
  wire [127:0] mem_7_io_memIO_rdata; // @[Top.scala 61:24]
  wire  block2_0 = riscvIns_block2_0;
  wire  _T = ~block2_0; // @[Top.scala 101:49]
  wire  _T_2 = ~riscvIns_io_instIO_ready; // @[Top.scala 257:37]
  wire  _T_3 = riscvIns_io_instIO_valid & _T_2; // @[Top.scala 257:34]
  wire  _T_4 = _T_3 ? axiIIO_io_axiIO_awvalid : axiDIO_io_axiIO_awvalid; // @[Top.scala 256:10]
  wire  DMABuzy_0 = dmaIns_DMABuzy_0;
  wire  _T_8 = _T_3 ? axiIIO_io_axiIO_wvalid : axiDIO_io_axiIO_wvalid; // @[Top.scala 256:10]
  wire  _T_12 = _T_3 ? axiIIO_io_axiIO_wlast : axiDIO_io_axiIO_wlast; // @[Top.scala 256:10]
  wire  _T_16 = _T_3 ? axiIIO_io_axiIO_bready : axiDIO_io_axiIO_bready; // @[Top.scala 256:10]
  wire  _T_20 = _T_3 ? axiIIO_io_axiIO_arvalid : axiDIO_io_axiIO_arvalid; // @[Top.scala 256:10]
  wire  _T_24 = _T_3 ? axiIIO_io_axiIO_rready : axiDIO_io_axiIO_rready; // @[Top.scala 256:10]
  wire [2:0] _T_32 = _T_3 ? axiIIO_io_axiIO_awsize : axiDIO_io_axiIO_awsize; // @[Top.scala 256:10]
  wire [31:0] _T_36 = _T_3 ? axiIIO_io_axiIO_awaddr : axiDIO_io_axiIO_awaddr; // @[Top.scala 256:10]
  wire [31:0] _T_40 = _T_3 ? axiIIO_io_axiIO_araddr : axiDIO_io_axiIO_araddr; // @[Top.scala 256:10]
  wire [63:0] _T_52 = _T_3 ? axiIIO_io_axiIO_wdata : axiDIO_io_axiIO_wdata; // @[Top.scala 256:10]
  wire [7:0] _T_60 = _T_3 ? axiIIO_io_axiIO_wstrb : axiDIO_io_axiIO_wstrb; // @[Top.scala 256:10]
  wire [7:0] _T_64 = _T_3 ? axiIIO_io_axiIO_arlen : axiDIO_io_axiIO_arlen; // @[Top.scala 256:10]
  wire [2:0] _T_68 = _T_3 ? axiIIO_io_axiIO_arsize : axiDIO_io_axiIO_arsize; // @[Top.scala 256:10]
  wire [1:0] _T_72 = _T_3 ? axiIIO_io_axiIO_arburst : axiDIO_io_axiIO_arburst; // @[Top.scala 256:10]
  wire  _T_77 = _T_3 | DMABuzy_0; // @[Top.scala 265:83]
  DMACtrl dmaIns ( // @[Top.scala 33:22]
    .clock(dmaIns_clock),
    .reset(dmaIns_reset),
    .io_dataIn_awready(dmaIns_io_dataIn_awready),
    .io_dataIn_awvalid(dmaIns_io_dataIn_awvalid),
    .io_dataIn_awaddr(dmaIns_io_dataIn_awaddr),
    .io_dataIn_awlen(dmaIns_io_dataIn_awlen),
    .io_dataIn_wready(dmaIns_io_dataIn_wready),
    .io_dataIn_wvalid(dmaIns_io_dataIn_wvalid),
    .io_dataIn_wdata(dmaIns_io_dataIn_wdata),
    .io_dataIn_wlast(dmaIns_io_dataIn_wlast),
    .io_dataIn_bready(dmaIns_io_dataIn_bready),
    .io_dataIn_bvalid(dmaIns_io_dataIn_bvalid),
    .io_dataIn_arready(dmaIns_io_dataIn_arready),
    .io_dataIn_arvalid(dmaIns_io_dataIn_arvalid),
    .io_dataIn_araddr(dmaIns_io_dataIn_araddr),
    .io_dataIn_arlen(dmaIns_io_dataIn_arlen),
    .io_dataIn_rready(dmaIns_io_dataIn_rready),
    .io_dataIn_rvalid(dmaIns_io_dataIn_rvalid),
    .io_dataIn_rdata(dmaIns_io_dataIn_rdata),
    .io_dataIn_rlast(dmaIns_io_dataIn_rlast),
    .io_dataOutMMIO_valid(dmaIns_io_dataOutMMIO_valid),
    .io_dataOutMMIO_ready(dmaIns_io_dataOutMMIO_ready),
    .io_dataOutMMIO_data_read(dmaIns_io_dataOutMMIO_data_read),
    .io_dataOutMMIO_data_write(dmaIns_io_dataOutMMIO_data_write),
    .io_dataOutMMIO_wen(dmaIns_io_dataOutMMIO_wen),
    .io_dataOutMMIO_addr(dmaIns_io_dataOutMMIO_addr),
    .dmaEn_0(dmaIns_dmaEn_0),
    .dmaEnWR_0(dmaIns_dmaEnWR_0),
    .block3_0(dmaIns_block3_0),
    .dmaCtrl_0(dmaIns_dmaCtrl_0),
    .block2_0(dmaIns_block2_0),
    .blockDMA_0(dmaIns_blockDMA_0),
    .DMABuzy_0(dmaIns_DMABuzy_0)
  );
  CGRAFullMask cgraIns ( // @[Top.scala 34:23]
    .clock(cgraIns_clock),
    .reset(cgraIns_reset),
    .io_CGRAIO_valid(cgraIns_io_CGRAIO_valid),
    .io_CGRAIO_ready(cgraIns_io_CGRAIO_ready),
    .io_CGRAIO_data_read(cgraIns_io_CGRAIO_data_read),
    .io_CGRAIO_data_write(cgraIns_io_CGRAIO_data_write),
    .io_CGRAIO_wen(cgraIns_io_CGRAIO_wen),
    .io_CGRAIO_addr(cgraIns_io_CGRAIO_addr),
    .io_outputs_0(cgraIns_io_outputs_0),
    .io_outputs_1(cgraIns_io_outputs_1),
    .io_outputs_2(cgraIns_io_outputs_2),
    .io_outputs_3(cgraIns_io_outputs_3),
    .io_outputs_4(cgraIns_io_outputs_4),
    .io_outputs_5(cgraIns_io_outputs_5),
    .io_outputs_6(cgraIns_io_outputs_6),
    .io_outputs_7(cgraIns_io_outputs_7),
    .io_outputs_8(cgraIns_io_outputs_8),
    .io_outputs_9(cgraIns_io_outputs_9),
    .io_outputs_10(cgraIns_io_outputs_10),
    .io_outputs_11(cgraIns_io_outputs_11),
    .io_outputs_12(cgraIns_io_outputs_12),
    .io_outputs_13(cgraIns_io_outputs_13),
    .io_outputs_14(cgraIns_io_outputs_14),
    .io_outputs_15(cgraIns_io_outputs_15),
    ._T_100_0(cgraIns__T_100_0),
    .dmaCtrl(cgraIns_dmaCtrl)
  );
  riscv riscvIns ( // @[Top.scala 35:24]
    .clock(riscvIns_clock),
    .reset(riscvIns_reset),
    .io_instIO_valid(riscvIns_io_instIO_valid),
    .io_instIO_ready(riscvIns_io_instIO_ready),
    .io_instIO_data_read(riscvIns_io_instIO_data_read),
    .io_instIO_addr(riscvIns_io_instIO_addr),
    .io_dataIO_valid(riscvIns_io_dataIO_valid),
    .io_dataIO_ready(riscvIns_io_dataIO_ready),
    .io_dataIO_data_read(riscvIns_io_dataIO_data_read),
    .io_dataIO_data_write(riscvIns_io_dataIO_data_write),
    .io_dataIO_wen(riscvIns_io_dataIO_wen),
    .io_dataIO_addr(riscvIns_io_dataIO_addr),
    .io_dataIO_rsize(riscvIns_io_dataIO_rsize),
    .io_dataIO_mask(riscvIns_io_dataIO_mask),
    ._T_99_0(riscvIns__T_99_0),
    .intrTimeCnt_0(riscvIns_intrTimeCnt_0),
    ._T_100_0(riscvIns__T_100_0),
    .startTimeCnt(riscvIns_startTimeCnt),
    .block3_0(riscvIns_block3_0),
    .dmaCtrl(riscvIns_dmaCtrl),
    .block2_0(riscvIns_block2_0),
    .blockDMA_0(riscvIns_blockDMA_0),
    .fencei_0(riscvIns_fencei_0)
  );
  Icache iCache ( // @[Top.scala 36:22]
    .clock(iCache_clock),
    .reset(iCache_reset),
    .io_cacheOut_ar_valid_o(iCache_io_cacheOut_ar_valid_o),
    .io_cacheOut_ar_addr_o(iCache_io_cacheOut_ar_addr_o),
    .io_cacheOut_ar_len_o(iCache_io_cacheOut_ar_len_o),
    .io_cacheOut_r_valid_i(iCache_io_cacheOut_r_valid_i),
    .io_cacheOut_r_data_i(iCache_io_cacheOut_r_data_i),
    .io_cacheOut_r_last_i(iCache_io_cacheOut_r_last_i),
    .io_cacheOut_w_addr_o(iCache_io_cacheOut_w_addr_o),
    .io_cacheIn_valid(iCache_io_cacheIn_valid),
    .io_cacheIn_ready(iCache_io_cacheIn_ready),
    .io_cacheIn_data_read(iCache_io_cacheIn_data_read),
    .io_cacheIn_addr(iCache_io_cacheIn_addr),
    .io_SRAMIO_0_cen(iCache_io_SRAMIO_0_cen),
    .io_SRAMIO_0_wen(iCache_io_SRAMIO_0_wen),
    .io_SRAMIO_0_wdata(iCache_io_SRAMIO_0_wdata),
    .io_SRAMIO_0_addr(iCache_io_SRAMIO_0_addr),
    .io_SRAMIO_0_wmask(iCache_io_SRAMIO_0_wmask),
    .io_SRAMIO_0_rdata(iCache_io_SRAMIO_0_rdata),
    .io_SRAMIO_1_cen(iCache_io_SRAMIO_1_cen),
    .io_SRAMIO_1_wen(iCache_io_SRAMIO_1_wen),
    .io_SRAMIO_1_wdata(iCache_io_SRAMIO_1_wdata),
    .io_SRAMIO_1_addr(iCache_io_SRAMIO_1_addr),
    .io_SRAMIO_1_wmask(iCache_io_SRAMIO_1_wmask),
    .io_SRAMIO_1_rdata(iCache_io_SRAMIO_1_rdata),
    .io_SRAMIO_2_cen(iCache_io_SRAMIO_2_cen),
    .io_SRAMIO_2_wen(iCache_io_SRAMIO_2_wen),
    .io_SRAMIO_2_wdata(iCache_io_SRAMIO_2_wdata),
    .io_SRAMIO_2_addr(iCache_io_SRAMIO_2_addr),
    .io_SRAMIO_2_wmask(iCache_io_SRAMIO_2_wmask),
    .io_SRAMIO_2_rdata(iCache_io_SRAMIO_2_rdata),
    .io_SRAMIO_3_cen(iCache_io_SRAMIO_3_cen),
    .io_SRAMIO_3_wen(iCache_io_SRAMIO_3_wen),
    .io_SRAMIO_3_wdata(iCache_io_SRAMIO_3_wdata),
    .io_SRAMIO_3_addr(iCache_io_SRAMIO_3_addr),
    .io_SRAMIO_3_wmask(iCache_io_SRAMIO_3_wmask),
    .io_SRAMIO_3_rdata(iCache_io_SRAMIO_3_rdata),
    .io_block(iCache_io_block),
    .updataICache(iCache_updataICache)
  );
  AXICache axiIIO ( // @[Top.scala 38:22]
    .clock(axiIIO_clock),
    .reset(axiIIO_reset),
    .io_axiIO_awready(axiIIO_io_axiIO_awready),
    .io_axiIO_awvalid(axiIIO_io_axiIO_awvalid),
    .io_axiIO_awaddr(axiIIO_io_axiIO_awaddr),
    .io_axiIO_awsize(axiIIO_io_axiIO_awsize),
    .io_axiIO_wready(axiIIO_io_axiIO_wready),
    .io_axiIO_wvalid(axiIIO_io_axiIO_wvalid),
    .io_axiIO_wdata(axiIIO_io_axiIO_wdata),
    .io_axiIO_wstrb(axiIIO_io_axiIO_wstrb),
    .io_axiIO_wlast(axiIIO_io_axiIO_wlast),
    .io_axiIO_bready(axiIIO_io_axiIO_bready),
    .io_axiIO_bvalid(axiIIO_io_axiIO_bvalid),
    .io_axiIO_arready(axiIIO_io_axiIO_arready),
    .io_axiIO_arvalid(axiIIO_io_axiIO_arvalid),
    .io_axiIO_araddr(axiIIO_io_axiIO_araddr),
    .io_axiIO_arlen(axiIIO_io_axiIO_arlen),
    .io_axiIO_arsize(axiIIO_io_axiIO_arsize),
    .io_axiIO_arburst(axiIIO_io_axiIO_arburst),
    .io_axiIO_rready(axiIIO_io_axiIO_rready),
    .io_axiIO_rvalid(axiIIO_io_axiIO_rvalid),
    .io_axiIO_rdata(axiIIO_io_axiIO_rdata),
    .io_axiIO_rlast(axiIIO_io_axiIO_rlast),
    .io_cache_ar_valid_o(axiIIO_io_cache_ar_valid_o),
    .io_cache_ar_addr_o(axiIIO_io_cache_ar_addr_o),
    .io_cache_ar_len_o(axiIIO_io_cache_ar_len_o),
    .io_cache_r_valid_i(axiIIO_io_cache_r_valid_i),
    .io_cache_r_data_i(axiIIO_io_cache_r_data_i),
    .io_cache_r_last_i(axiIIO_io_cache_r_last_i),
    .io_cache_w_valid_o(axiIIO_io_cache_w_valid_o),
    .io_cache_w_ready_i(axiIIO_io_cache_w_ready_i),
    .io_cache_w_data_o(axiIIO_io_cache_w_data_o),
    .io_cache_w_addr_o(axiIIO_io_cache_w_addr_o),
    .io_cache_w_mask_o(axiIIO_io_cache_w_mask_o),
    .io_cache_wsize(axiIIO_io_cache_wsize)
  );
  arbTop dArbIns ( // @[Top.scala 41:23]
    .io_arbIn_valid(dArbIns_io_arbIn_valid),
    .io_arbIn_ready(dArbIns_io_arbIn_ready),
    .io_arbIn_data_read(dArbIns_io_arbIn_data_read),
    .io_arbIn_data_write(dArbIns_io_arbIn_data_write),
    .io_arbIn_wen(dArbIns_io_arbIn_wen),
    .io_arbIn_addr(dArbIns_io_arbIn_addr),
    .io_arbIn_rsize(dArbIns_io_arbIn_rsize),
    .io_arbIn_mask(dArbIns_io_arbIn_mask),
    .io_arbMMIO_valid(dArbIns_io_arbMMIO_valid),
    .io_arbMMIO_ready(dArbIns_io_arbMMIO_ready),
    .io_arbMMIO_data_read(dArbIns_io_arbMMIO_data_read),
    .io_arbMMIO_data_write(dArbIns_io_arbMMIO_data_write),
    .io_arbMMIO_wen(dArbIns_io_arbMMIO_wen),
    .io_arbMMIO_addr(dArbIns_io_arbMMIO_addr),
    .io_arbMMIO_rsize(dArbIns_io_arbMMIO_rsize),
    .io_arbMMIO_mask(dArbIns_io_arbMMIO_mask),
    .io_arbClint_valid(dArbIns_io_arbClint_valid),
    .io_arbClint_data_read(dArbIns_io_arbClint_data_read),
    .io_arbClint_data_write(dArbIns_io_arbClint_data_write),
    .io_arbClint_wen(dArbIns_io_arbClint_wen),
    .io_arbClint_addr(dArbIns_io_arbClint_addr),
    .io_arbDCache_valid(dArbIns_io_arbDCache_valid),
    .io_arbDCache_ready(dArbIns_io_arbDCache_ready),
    .io_arbDCache_data_read(dArbIns_io_arbDCache_data_read),
    .io_arbDCache_data_write(dArbIns_io_arbDCache_data_write),
    .io_arbDCache_wen(dArbIns_io_arbDCache_wen),
    .io_arbDCache_addr(dArbIns_io_arbDCache_addr),
    .io_arbDCache_rsize(dArbIns_io_arbDCache_rsize),
    .io_arbDCache_mask(dArbIns_io_arbDCache_mask),
    .io_arbCgra_valid(dArbIns_io_arbCgra_valid),
    .io_arbCgra_ready(dArbIns_io_arbCgra_ready),
    .io_arbCgra_data_read(dArbIns_io_arbCgra_data_read),
    .io_arbCgra_data_write(dArbIns_io_arbCgra_data_write),
    .io_arbCgra_wen(dArbIns_io_arbCgra_wen),
    .io_arbCgra_addr(dArbIns_io_arbCgra_addr)
  );
  mmioCache mmioDCache ( // @[Top.scala 42:26]
    .io_mmioIn_valid(mmioDCache_io_mmioIn_valid),
    .io_mmioIn_ready(mmioDCache_io_mmioIn_ready),
    .io_mmioIn_data_read(mmioDCache_io_mmioIn_data_read),
    .io_mmioIn_data_write(mmioDCache_io_mmioIn_data_write),
    .io_mmioIn_wen(mmioDCache_io_mmioIn_wen),
    .io_mmioIn_addr(mmioDCache_io_mmioIn_addr),
    .io_mmioOut_valid(mmioDCache_io_mmioOut_valid),
    .io_mmioOut_ready(mmioDCache_io_mmioOut_ready),
    .io_mmioOut_data_read(mmioDCache_io_mmioOut_data_read),
    .io_mmioOut_data_write(mmioDCache_io_mmioOut_data_write),
    .io_mmioOut_wen(mmioDCache_io_mmioOut_wen),
    .io_mmioOut_addr(mmioDCache_io_mmioOut_addr)
  );
  Dcache dCache ( // @[Top.scala 43:22]
    .clock(dCache_clock),
    .reset(dCache_reset),
    .io_cacheOut_ar_valid_o(dCache_io_cacheOut_ar_valid_o),
    .io_cacheOut_ar_addr_o(dCache_io_cacheOut_ar_addr_o),
    .io_cacheOut_ar_len_o(dCache_io_cacheOut_ar_len_o),
    .io_cacheOut_r_valid_i(dCache_io_cacheOut_r_valid_i),
    .io_cacheOut_r_data_i(dCache_io_cacheOut_r_data_i),
    .io_cacheOut_r_last_i(dCache_io_cacheOut_r_last_i),
    .io_cacheOut_w_valid_o(dCache_io_cacheOut_w_valid_o),
    .io_cacheOut_w_ready_i(dCache_io_cacheOut_w_ready_i),
    .io_cacheOut_w_data_o(dCache_io_cacheOut_w_data_o),
    .io_cacheOut_w_addr_o(dCache_io_cacheOut_w_addr_o),
    .io_cacheOut_w_mask_o(dCache_io_cacheOut_w_mask_o),
    .io_cacheOut_wsize(dCache_io_cacheOut_wsize),
    .io_cacheIn_valid(dCache_io_cacheIn_valid),
    .io_cacheIn_ready(dCache_io_cacheIn_ready),
    .io_cacheIn_data_read(dCache_io_cacheIn_data_read),
    .io_cacheIn_data_write(dCache_io_cacheIn_data_write),
    .io_cacheIn_wen(dCache_io_cacheIn_wen),
    .io_cacheIn_addr(dCache_io_cacheIn_addr),
    .io_cacheIn_rsize(dCache_io_cacheIn_rsize),
    .io_cacheIn_mask(dCache_io_cacheIn_mask),
    .io_SRAMIO_0_cen(dCache_io_SRAMIO_0_cen),
    .io_SRAMIO_0_wen(dCache_io_SRAMIO_0_wen),
    .io_SRAMIO_0_wdata(dCache_io_SRAMIO_0_wdata),
    .io_SRAMIO_0_addr(dCache_io_SRAMIO_0_addr),
    .io_SRAMIO_0_wmask(dCache_io_SRAMIO_0_wmask),
    .io_SRAMIO_0_rdata(dCache_io_SRAMIO_0_rdata),
    .io_SRAMIO_1_cen(dCache_io_SRAMIO_1_cen),
    .io_SRAMIO_1_wen(dCache_io_SRAMIO_1_wen),
    .io_SRAMIO_1_wdata(dCache_io_SRAMIO_1_wdata),
    .io_SRAMIO_1_addr(dCache_io_SRAMIO_1_addr),
    .io_SRAMIO_1_wmask(dCache_io_SRAMIO_1_wmask),
    .io_SRAMIO_1_rdata(dCache_io_SRAMIO_1_rdata),
    .io_SRAMIO_2_cen(dCache_io_SRAMIO_2_cen),
    .io_SRAMIO_2_wen(dCache_io_SRAMIO_2_wen),
    .io_SRAMIO_2_wdata(dCache_io_SRAMIO_2_wdata),
    .io_SRAMIO_2_addr(dCache_io_SRAMIO_2_addr),
    .io_SRAMIO_2_wmask(dCache_io_SRAMIO_2_wmask),
    .io_SRAMIO_2_rdata(dCache_io_SRAMIO_2_rdata),
    .io_SRAMIO_3_cen(dCache_io_SRAMIO_3_cen),
    .io_SRAMIO_3_wen(dCache_io_SRAMIO_3_wen),
    .io_SRAMIO_3_wdata(dCache_io_SRAMIO_3_wdata),
    .io_SRAMIO_3_addr(dCache_io_SRAMIO_3_addr),
    .io_SRAMIO_3_wmask(dCache_io_SRAMIO_3_wmask),
    .io_SRAMIO_3_rdata(dCache_io_SRAMIO_3_rdata),
    .io_block(dCache_io_block),
    .updataICache(dCache_updataICache)
  );
  clint clintIns ( // @[Top.scala 44:25]
    .clock(clintIns_clock),
    .reset(clintIns_reset),
    .io_clintIO_valid(clintIns_io_clintIO_valid),
    .io_clintIO_data_read(clintIns_io_clintIO_data_read),
    .io_clintIO_data_write(clintIns_io_clintIO_data_write),
    .io_clintIO_wen(clintIns_io_clintIO_wen),
    .io_clintIO_addr(clintIns_io_clintIO_addr),
    .intrTimeCnt_0(clintIns_intrTimeCnt_0),
    .startTimeCnt_0(clintIns_startTimeCnt_0)
  );
  AXICache axiDIO ( // @[Top.scala 53:22]
    .clock(axiDIO_clock),
    .reset(axiDIO_reset),
    .io_axiIO_awready(axiDIO_io_axiIO_awready),
    .io_axiIO_awvalid(axiDIO_io_axiIO_awvalid),
    .io_axiIO_awaddr(axiDIO_io_axiIO_awaddr),
    .io_axiIO_awsize(axiDIO_io_axiIO_awsize),
    .io_axiIO_wready(axiDIO_io_axiIO_wready),
    .io_axiIO_wvalid(axiDIO_io_axiIO_wvalid),
    .io_axiIO_wdata(axiDIO_io_axiIO_wdata),
    .io_axiIO_wstrb(axiDIO_io_axiIO_wstrb),
    .io_axiIO_wlast(axiDIO_io_axiIO_wlast),
    .io_axiIO_bready(axiDIO_io_axiIO_bready),
    .io_axiIO_bvalid(axiDIO_io_axiIO_bvalid),
    .io_axiIO_arready(axiDIO_io_axiIO_arready),
    .io_axiIO_arvalid(axiDIO_io_axiIO_arvalid),
    .io_axiIO_araddr(axiDIO_io_axiIO_araddr),
    .io_axiIO_arlen(axiDIO_io_axiIO_arlen),
    .io_axiIO_arsize(axiDIO_io_axiIO_arsize),
    .io_axiIO_arburst(axiDIO_io_axiIO_arburst),
    .io_axiIO_rready(axiDIO_io_axiIO_rready),
    .io_axiIO_rvalid(axiDIO_io_axiIO_rvalid),
    .io_axiIO_rdata(axiDIO_io_axiIO_rdata),
    .io_axiIO_rlast(axiDIO_io_axiIO_rlast),
    .io_cache_ar_valid_o(axiDIO_io_cache_ar_valid_o),
    .io_cache_ar_addr_o(axiDIO_io_cache_ar_addr_o),
    .io_cache_ar_len_o(axiDIO_io_cache_ar_len_o),
    .io_cache_r_valid_i(axiDIO_io_cache_r_valid_i),
    .io_cache_r_data_i(axiDIO_io_cache_r_data_i),
    .io_cache_r_last_i(axiDIO_io_cache_r_last_i),
    .io_cache_w_valid_o(axiDIO_io_cache_w_valid_o),
    .io_cache_w_ready_i(axiDIO_io_cache_w_ready_i),
    .io_cache_w_data_o(axiDIO_io_cache_w_data_o),
    .io_cache_w_addr_o(axiDIO_io_cache_w_addr_o),
    .io_cache_w_mask_o(axiDIO_io_cache_w_mask_o),
    .io_cache_wsize(axiDIO_io_cache_wsize)
  );
  mem mem ( // @[Top.scala 60:24]
    .clock(mem_clock),
    .io_memIO_cen(mem_io_memIO_cen),
    .io_memIO_wen(mem_io_memIO_wen),
    .io_memIO_wdata(mem_io_memIO_wdata),
    .io_memIO_addr(mem_io_memIO_addr),
    .io_memIO_wmask(mem_io_memIO_wmask),
    .io_memIO_rdata(mem_io_memIO_rdata)
  );
  mem mem_1 ( // @[Top.scala 61:24]
    .clock(mem_1_clock),
    .io_memIO_cen(mem_1_io_memIO_cen),
    .io_memIO_wen(mem_1_io_memIO_wen),
    .io_memIO_wdata(mem_1_io_memIO_wdata),
    .io_memIO_addr(mem_1_io_memIO_addr),
    .io_memIO_wmask(mem_1_io_memIO_wmask),
    .io_memIO_rdata(mem_1_io_memIO_rdata)
  );
  mem mem_2 ( // @[Top.scala 60:24]
    .clock(mem_2_clock),
    .io_memIO_cen(mem_2_io_memIO_cen),
    .io_memIO_wen(mem_2_io_memIO_wen),
    .io_memIO_wdata(mem_2_io_memIO_wdata),
    .io_memIO_addr(mem_2_io_memIO_addr),
    .io_memIO_wmask(mem_2_io_memIO_wmask),
    .io_memIO_rdata(mem_2_io_memIO_rdata)
  );
  mem mem_3 ( // @[Top.scala 61:24]
    .clock(mem_3_clock),
    .io_memIO_cen(mem_3_io_memIO_cen),
    .io_memIO_wen(mem_3_io_memIO_wen),
    .io_memIO_wdata(mem_3_io_memIO_wdata),
    .io_memIO_addr(mem_3_io_memIO_addr),
    .io_memIO_wmask(mem_3_io_memIO_wmask),
    .io_memIO_rdata(mem_3_io_memIO_rdata)
  );
  mem mem_4 ( // @[Top.scala 60:24]
    .clock(mem_4_clock),
    .io_memIO_cen(mem_4_io_memIO_cen),
    .io_memIO_wen(mem_4_io_memIO_wen),
    .io_memIO_wdata(mem_4_io_memIO_wdata),
    .io_memIO_addr(mem_4_io_memIO_addr),
    .io_memIO_wmask(mem_4_io_memIO_wmask),
    .io_memIO_rdata(mem_4_io_memIO_rdata)
  );
  mem mem_5 ( // @[Top.scala 61:24]
    .clock(mem_5_clock),
    .io_memIO_cen(mem_5_io_memIO_cen),
    .io_memIO_wen(mem_5_io_memIO_wen),
    .io_memIO_wdata(mem_5_io_memIO_wdata),
    .io_memIO_addr(mem_5_io_memIO_addr),
    .io_memIO_wmask(mem_5_io_memIO_wmask),
    .io_memIO_rdata(mem_5_io_memIO_rdata)
  );
  mem mem_6 ( // @[Top.scala 60:24]
    .clock(mem_6_clock),
    .io_memIO_cen(mem_6_io_memIO_cen),
    .io_memIO_wen(mem_6_io_memIO_wen),
    .io_memIO_wdata(mem_6_io_memIO_wdata),
    .io_memIO_addr(mem_6_io_memIO_addr),
    .io_memIO_wmask(mem_6_io_memIO_wmask),
    .io_memIO_rdata(mem_6_io_memIO_rdata)
  );
  mem mem_7 ( // @[Top.scala 61:24]
    .clock(mem_7_clock),
    .io_memIO_cen(mem_7_io_memIO_cen),
    .io_memIO_wen(mem_7_io_memIO_wen),
    .io_memIO_wdata(mem_7_io_memIO_wdata),
    .io_memIO_addr(mem_7_io_memIO_addr),
    .io_memIO_wmask(mem_7_io_memIO_wmask),
    .io_memIO_rdata(mem_7_io_memIO_rdata)
  );
  assign io_dmaster_awvalid = DMABuzy_0 ? dmaIns_io_dataIn_awvalid : _T_4; // @[Top.scala 253:23]
  assign io_dmaster_awid = 4'h0; // @[Top.scala 253:23]
  assign io_dmaster_awaddr = DMABuzy_0 ? dmaIns_io_dataIn_awaddr : _T_36; // @[Top.scala 253:23]
  assign io_dmaster_awlen = DMABuzy_0 ? dmaIns_io_dataIn_awlen : 8'h0; // @[Top.scala 253:23]
  assign io_dmaster_awsize = DMABuzy_0 ? 3'h3 : _T_32; // @[Top.scala 253:23]
  assign io_dmaster_awburst = 2'h1; // @[Top.scala 253:23]
  assign io_dmaster_wvalid = DMABuzy_0 ? dmaIns_io_dataIn_wvalid : _T_8; // @[Top.scala 253:23]
  assign io_dmaster_wdata = DMABuzy_0 ? dmaIns_io_dataIn_wdata : _T_52; // @[Top.scala 253:23]
  assign io_dmaster_wstrb = DMABuzy_0 ? 8'hff : _T_60; // @[Top.scala 253:23]
  assign io_dmaster_wlast = DMABuzy_0 ? dmaIns_io_dataIn_wlast : _T_12; // @[Top.scala 253:23]
  assign io_dmaster_bready = DMABuzy_0 ? dmaIns_io_dataIn_bready : _T_16; // @[Top.scala 253:23]
  assign io_dmaster_arvalid = DMABuzy_0 ? dmaIns_io_dataIn_arvalid : _T_20; // @[Top.scala 253:23]
  assign io_dmaster_arid = 4'h0; // @[Top.scala 253:23]
  assign io_dmaster_araddr = DMABuzy_0 ? dmaIns_io_dataIn_araddr : _T_40; // @[Top.scala 253:23]
  assign io_dmaster_arlen = DMABuzy_0 ? dmaIns_io_dataIn_arlen : _T_64; // @[Top.scala 253:23]
  assign io_dmaster_arsize = DMABuzy_0 ? 3'h3 : _T_68; // @[Top.scala 253:23]
  assign io_dmaster_arburst = DMABuzy_0 ? 2'h1 : _T_72; // @[Top.scala 253:23]
  assign io_dmaster_rready = DMABuzy_0 ? dmaIns_io_dataIn_rready : _T_24; // @[Top.scala 253:23]
  assign io_outputs_0 = cgraIns_io_outputs_0; // @[Top.scala 45:14]
  assign io_outputs_1 = cgraIns_io_outputs_1; // @[Top.scala 45:14]
  assign io_outputs_2 = cgraIns_io_outputs_2; // @[Top.scala 45:14]
  assign io_outputs_3 = cgraIns_io_outputs_3; // @[Top.scala 45:14]
  assign io_outputs_4 = cgraIns_io_outputs_4; // @[Top.scala 45:14]
  assign io_outputs_5 = cgraIns_io_outputs_5; // @[Top.scala 45:14]
  assign io_outputs_6 = cgraIns_io_outputs_6; // @[Top.scala 45:14]
  assign io_outputs_7 = cgraIns_io_outputs_7; // @[Top.scala 45:14]
  assign io_outputs_8 = cgraIns_io_outputs_8; // @[Top.scala 45:14]
  assign io_outputs_9 = cgraIns_io_outputs_9; // @[Top.scala 45:14]
  assign io_outputs_10 = cgraIns_io_outputs_10; // @[Top.scala 45:14]
  assign io_outputs_11 = cgraIns_io_outputs_11; // @[Top.scala 45:14]
  assign io_outputs_12 = cgraIns_io_outputs_12; // @[Top.scala 45:14]
  assign io_outputs_13 = cgraIns_io_outputs_13; // @[Top.scala 45:14]
  assign io_outputs_14 = cgraIns_io_outputs_14; // @[Top.scala 45:14]
  assign io_outputs_15 = cgraIns_io_outputs_15; // @[Top.scala 45:14]
  assign io_mmio_valid = dArbIns_io_arbMMIO_valid & _T; // @[Top.scala 50:21 Top.scala 101:17]
  assign io_mmio_data_write = dArbIns_io_arbMMIO_data_write; // @[Top.scala 50:21]
  assign io_mmio_wen = dArbIns_io_arbMMIO_wen; // @[Top.scala 50:21]
  assign io_mmio_addr = dArbIns_io_arbMMIO_addr; // @[Top.scala 50:21]
  assign io_mmio_rsize = dArbIns_io_arbMMIO_rsize; // @[Top.scala 50:21]
  assign io_mmio_mask = dArbIns_io_arbMMIO_mask; // @[Top.scala 50:21]
  assign dmaIns_clock = clock;
  assign dmaIns_reset = reset;
  assign dmaIns_io_dataIn_awready = io_dmaster_awready; // @[Top.scala 263:21]
  assign dmaIns_io_dataIn_wready = io_dmaster_wready; // @[Top.scala 263:21]
  assign dmaIns_io_dataIn_bvalid = io_dmaster_bvalid; // @[Top.scala 263:21]
  assign dmaIns_io_dataIn_arready = io_dmaster_arready; // @[Top.scala 263:21]
  assign dmaIns_io_dataIn_rvalid = io_dmaster_rvalid; // @[Top.scala 263:21]
  assign dmaIns_io_dataIn_rdata = io_dmaster_rdata; // @[Top.scala 263:21]
  assign dmaIns_io_dataIn_rlast = io_dmaster_rlast; // @[Top.scala 263:21]
  assign dmaIns_io_dataOutMMIO_ready = cgraIns_io_CGRAIO_ready; // @[Top.scala 318:22]
  assign dmaIns_io_dataOutMMIO_data_read = cgraIns_io_CGRAIO_data_read; // @[Top.scala 318:22]
  assign dmaIns_dmaEn_0 = riscvIns__T_99_0;
  assign dmaIns_dmaEnWR_0 = riscvIns__T_100_0;
  assign dmaIns_block3_0 = riscvIns_block3_0;
  assign dmaIns_dmaCtrl_0 = riscvIns_dmaCtrl;
  assign dmaIns_block2_0 = riscvIns_block2_0;
  assign cgraIns_clock = clock;
  assign cgraIns_reset = reset;
  assign cgraIns_io_CGRAIO_valid = DMABuzy_0 ? dmaIns_io_dataOutMMIO_valid : mmioDCache_io_mmioOut_valid; // @[Top.scala 311:22]
  assign cgraIns_io_CGRAIO_data_write = DMABuzy_0 ? dmaIns_io_dataOutMMIO_data_write : mmioDCache_io_mmioOut_data_write; // @[Top.scala 311:22]
  assign cgraIns_io_CGRAIO_wen = DMABuzy_0 ? dmaIns_io_dataOutMMIO_wen : mmioDCache_io_mmioOut_wen; // @[Top.scala 311:22]
  assign cgraIns_io_CGRAIO_addr = DMABuzy_0 ? dmaIns_io_dataOutMMIO_addr : mmioDCache_io_mmioOut_addr; // @[Top.scala 311:22]
  assign cgraIns__T_100_0 = riscvIns__T_100_0;
  assign cgraIns_dmaCtrl = riscvIns_dmaCtrl;
  assign riscvIns_clock = clock;
  assign riscvIns_reset = reset;
  assign riscvIns_io_instIO_ready = iCache_io_cacheIn_ready; // @[Top.scala 37:22]
  assign riscvIns_io_instIO_data_read = iCache_io_cacheIn_data_read; // @[Top.scala 37:22]
  assign riscvIns_io_dataIO_ready = dArbIns_io_arbIn_ready; // @[Top.scala 46:21]
  assign riscvIns_io_dataIO_data_read = dArbIns_io_arbIn_data_read; // @[Top.scala 46:21]
  assign riscvIns_intrTimeCnt_0 = clintIns_intrTimeCnt_0;
  assign riscvIns_blockDMA_0 = dmaIns_blockDMA_0;
  assign iCache_clock = clock;
  assign iCache_reset = reset;
  assign iCache_io_cacheOut_r_valid_i = axiIIO_io_cache_r_valid_i; // @[Top.scala 39:19]
  assign iCache_io_cacheOut_r_data_i = axiIIO_io_cache_r_data_i; // @[Top.scala 39:19]
  assign iCache_io_cacheOut_r_last_i = axiIIO_io_cache_r_last_i; // @[Top.scala 39:19]
  assign iCache_io_cacheIn_valid = riscvIns_io_instIO_valid; // @[Top.scala 37:22]
  assign iCache_io_cacheIn_addr = riscvIns_io_instIO_addr; // @[Top.scala 37:22]
  assign iCache_io_SRAMIO_0_rdata = mem_io_memIO_rdata; // @[Top.scala 62:20]
  assign iCache_io_SRAMIO_1_rdata = mem_2_io_memIO_rdata; // @[Top.scala 62:20]
  assign iCache_io_SRAMIO_2_rdata = mem_4_io_memIO_rdata; // @[Top.scala 62:20]
  assign iCache_io_SRAMIO_3_rdata = mem_6_io_memIO_rdata; // @[Top.scala 62:20]
  assign iCache_io_block = riscvIns_block3_0; // @[Top.scala 98:21]
  assign iCache_updataICache = riscvIns_fencei_0;
  assign axiIIO_clock = clock;
  assign axiIIO_reset = reset;
  assign axiIIO_io_axiIO_awready = DMABuzy_0 ? 1'h0 : io_dmaster_awready; // @[Top.scala 264:24]
  assign axiIIO_io_axiIO_wready = DMABuzy_0 ? 1'h0 : io_dmaster_wready; // @[Top.scala 264:24]
  assign axiIIO_io_axiIO_bvalid = DMABuzy_0 ? 1'h0 : io_dmaster_bvalid; // @[Top.scala 264:24]
  assign axiIIO_io_axiIO_arready = DMABuzy_0 ? 1'h0 : io_dmaster_arready; // @[Top.scala 264:24]
  assign axiIIO_io_axiIO_rvalid = DMABuzy_0 ? 1'h0 : io_dmaster_rvalid; // @[Top.scala 264:24]
  assign axiIIO_io_axiIO_rdata = DMABuzy_0 ? 64'h0 : io_dmaster_rdata; // @[Top.scala 264:24]
  assign axiIIO_io_axiIO_rlast = DMABuzy_0 ? 1'h0 : io_dmaster_rlast; // @[Top.scala 264:24]
  assign axiIIO_io_cache_ar_valid_o = iCache_io_cacheOut_ar_valid_o; // @[Top.scala 39:19]
  assign axiIIO_io_cache_ar_addr_o = iCache_io_cacheOut_ar_addr_o; // @[Top.scala 39:19]
  assign axiIIO_io_cache_ar_len_o = iCache_io_cacheOut_ar_len_o; // @[Top.scala 39:19]
  assign axiIIO_io_cache_w_valid_o = 1'h0; // @[Top.scala 39:19]
  assign axiIIO_io_cache_w_data_o = 64'h0; // @[Top.scala 39:19]
  assign axiIIO_io_cache_w_addr_o = iCache_io_cacheOut_w_addr_o; // @[Top.scala 39:19]
  assign axiIIO_io_cache_w_mask_o = 8'h0; // @[Top.scala 39:19]
  assign axiIIO_io_cache_wsize = 2'h2; // @[Top.scala 39:19]
  assign dArbIns_io_arbIn_valid = riscvIns_io_dataIO_valid; // @[Top.scala 46:21]
  assign dArbIns_io_arbIn_data_write = riscvIns_io_dataIO_data_write; // @[Top.scala 46:21]
  assign dArbIns_io_arbIn_wen = riscvIns_io_dataIO_wen; // @[Top.scala 46:21]
  assign dArbIns_io_arbIn_addr = riscvIns_io_dataIO_addr; // @[Top.scala 46:21]
  assign dArbIns_io_arbIn_rsize = riscvIns_io_dataIO_rsize; // @[Top.scala 46:21]
  assign dArbIns_io_arbIn_mask = riscvIns_io_dataIO_mask; // @[Top.scala 46:21]
  assign dArbIns_io_arbMMIO_ready = io_mmio_ready; // @[Top.scala 50:21]
  assign dArbIns_io_arbMMIO_data_read = io_mmio_data_read; // @[Top.scala 50:21]
  assign dArbIns_io_arbClint_data_read = clintIns_io_clintIO_data_read; // @[Top.scala 49:22]
  assign dArbIns_io_arbDCache_ready = dCache_io_cacheIn_ready; // @[Top.scala 48:24]
  assign dArbIns_io_arbDCache_data_read = dCache_io_cacheIn_data_read; // @[Top.scala 48:24]
  assign dArbIns_io_arbCgra_ready = mmioDCache_io_mmioIn_ready; // @[Top.scala 47:21]
  assign dArbIns_io_arbCgra_data_read = mmioDCache_io_mmioIn_data_read; // @[Top.scala 47:21]
  assign mmioDCache_io_mmioIn_valid = dArbIns_io_arbCgra_valid; // @[Top.scala 47:21]
  assign mmioDCache_io_mmioIn_data_write = dArbIns_io_arbCgra_data_write; // @[Top.scala 47:21]
  assign mmioDCache_io_mmioIn_wen = dArbIns_io_arbCgra_wen; // @[Top.scala 47:21]
  assign mmioDCache_io_mmioIn_addr = dArbIns_io_arbCgra_addr; // @[Top.scala 47:21]
  assign mmioDCache_io_mmioOut_ready = cgraIns_io_CGRAIO_ready; // @[Top.scala 319:25]
  assign mmioDCache_io_mmioOut_data_read = cgraIns_io_CGRAIO_data_read; // @[Top.scala 319:25]
  assign dCache_clock = clock;
  assign dCache_reset = reset;
  assign dCache_io_cacheOut_r_valid_i = axiDIO_io_cache_r_valid_i; // @[Top.scala 55:18]
  assign dCache_io_cacheOut_r_data_i = axiDIO_io_cache_r_data_i; // @[Top.scala 55:18]
  assign dCache_io_cacheOut_r_last_i = axiDIO_io_cache_r_last_i; // @[Top.scala 55:18]
  assign dCache_io_cacheOut_w_ready_i = axiDIO_io_cache_w_ready_i; // @[Top.scala 55:18]
  assign dCache_io_cacheIn_valid = dArbIns_io_arbDCache_valid; // @[Top.scala 48:24]
  assign dCache_io_cacheIn_data_write = dArbIns_io_arbDCache_data_write; // @[Top.scala 48:24]
  assign dCache_io_cacheIn_wen = dArbIns_io_arbDCache_wen; // @[Top.scala 48:24]
  assign dCache_io_cacheIn_addr = dArbIns_io_arbDCache_addr; // @[Top.scala 48:24]
  assign dCache_io_cacheIn_rsize = dArbIns_io_arbDCache_rsize; // @[Top.scala 48:24]
  assign dCache_io_cacheIn_mask = dArbIns_io_arbDCache_mask; // @[Top.scala 48:24]
  assign dCache_io_SRAMIO_0_rdata = mem_1_io_memIO_rdata; // @[Top.scala 63:20]
  assign dCache_io_SRAMIO_1_rdata = mem_3_io_memIO_rdata; // @[Top.scala 63:20]
  assign dCache_io_SRAMIO_2_rdata = mem_5_io_memIO_rdata; // @[Top.scala 63:20]
  assign dCache_io_SRAMIO_3_rdata = mem_7_io_memIO_rdata; // @[Top.scala 63:20]
  assign dCache_io_block = riscvIns_block2_0; // @[Top.scala 100:19]
  assign dCache_updataICache = riscvIns_fencei_0;
  assign clintIns_clock = clock;
  assign clintIns_reset = reset;
  assign clintIns_io_clintIO_valid = dArbIns_io_arbClint_valid; // @[Top.scala 49:22]
  assign clintIns_io_clintIO_data_write = dArbIns_io_arbClint_data_write; // @[Top.scala 49:22]
  assign clintIns_io_clintIO_wen = dArbIns_io_arbClint_wen; // @[Top.scala 49:22]
  assign clintIns_io_clintIO_addr = dArbIns_io_arbClint_addr; // @[Top.scala 49:22]
  assign clintIns_startTimeCnt_0 = riscvIns_startTimeCnt;
  assign axiDIO_clock = clock;
  assign axiDIO_reset = reset;
  assign axiDIO_io_axiIO_awready = _T_77 ? 1'h0 : io_dmaster_awready; // @[Top.scala 265:21]
  assign axiDIO_io_axiIO_wready = _T_77 ? 1'h0 : io_dmaster_wready; // @[Top.scala 265:21]
  assign axiDIO_io_axiIO_bvalid = _T_77 ? 1'h0 : io_dmaster_bvalid; // @[Top.scala 265:21]
  assign axiDIO_io_axiIO_arready = _T_77 ? 1'h0 : io_dmaster_arready; // @[Top.scala 265:21]
  assign axiDIO_io_axiIO_rvalid = _T_77 ? 1'h0 : io_dmaster_rvalid; // @[Top.scala 265:21]
  assign axiDIO_io_axiIO_rdata = _T_77 ? 64'h0 : io_dmaster_rdata; // @[Top.scala 265:21]
  assign axiDIO_io_axiIO_rlast = _T_77 ? 1'h0 : io_dmaster_rlast; // @[Top.scala 265:21]
  assign axiDIO_io_cache_ar_valid_o = dCache_io_cacheOut_ar_valid_o; // @[Top.scala 55:18]
  assign axiDIO_io_cache_ar_addr_o = dCache_io_cacheOut_ar_addr_o; // @[Top.scala 55:18]
  assign axiDIO_io_cache_ar_len_o = dCache_io_cacheOut_ar_len_o; // @[Top.scala 55:18]
  assign axiDIO_io_cache_w_valid_o = dCache_io_cacheOut_w_valid_o; // @[Top.scala 55:18]
  assign axiDIO_io_cache_w_data_o = dCache_io_cacheOut_w_data_o; // @[Top.scala 55:18]
  assign axiDIO_io_cache_w_addr_o = dCache_io_cacheOut_w_addr_o; // @[Top.scala 55:18]
  assign axiDIO_io_cache_w_mask_o = dCache_io_cacheOut_w_mask_o; // @[Top.scala 55:18]
  assign axiDIO_io_cache_wsize = dCache_io_cacheOut_wsize; // @[Top.scala 55:18]
  assign mem_clock = clock;
  assign mem_io_memIO_cen = iCache_io_SRAMIO_0_cen; // @[Top.scala 62:20]
  assign mem_io_memIO_wen = iCache_io_SRAMIO_0_wen; // @[Top.scala 62:20]
  assign mem_io_memIO_wdata = iCache_io_SRAMIO_0_wdata; // @[Top.scala 62:20]
  assign mem_io_memIO_addr = iCache_io_SRAMIO_0_addr; // @[Top.scala 62:20]
  assign mem_io_memIO_wmask = iCache_io_SRAMIO_0_wmask; // @[Top.scala 62:20]
  assign mem_1_clock = clock;
  assign mem_1_io_memIO_cen = dCache_io_SRAMIO_0_cen; // @[Top.scala 63:20]
  assign mem_1_io_memIO_wen = dCache_io_SRAMIO_0_wen; // @[Top.scala 63:20]
  assign mem_1_io_memIO_wdata = dCache_io_SRAMIO_0_wdata; // @[Top.scala 63:20]
  assign mem_1_io_memIO_addr = dCache_io_SRAMIO_0_addr; // @[Top.scala 63:20]
  assign mem_1_io_memIO_wmask = dCache_io_SRAMIO_0_wmask; // @[Top.scala 63:20]
  assign mem_2_clock = clock;
  assign mem_2_io_memIO_cen = iCache_io_SRAMIO_1_cen; // @[Top.scala 62:20]
  assign mem_2_io_memIO_wen = iCache_io_SRAMIO_1_wen; // @[Top.scala 62:20]
  assign mem_2_io_memIO_wdata = iCache_io_SRAMIO_1_wdata; // @[Top.scala 62:20]
  assign mem_2_io_memIO_addr = iCache_io_SRAMIO_1_addr; // @[Top.scala 62:20]
  assign mem_2_io_memIO_wmask = iCache_io_SRAMIO_1_wmask; // @[Top.scala 62:20]
  assign mem_3_clock = clock;
  assign mem_3_io_memIO_cen = dCache_io_SRAMIO_1_cen; // @[Top.scala 63:20]
  assign mem_3_io_memIO_wen = dCache_io_SRAMIO_1_wen; // @[Top.scala 63:20]
  assign mem_3_io_memIO_wdata = dCache_io_SRAMIO_1_wdata; // @[Top.scala 63:20]
  assign mem_3_io_memIO_addr = dCache_io_SRAMIO_1_addr; // @[Top.scala 63:20]
  assign mem_3_io_memIO_wmask = dCache_io_SRAMIO_1_wmask; // @[Top.scala 63:20]
  assign mem_4_clock = clock;
  assign mem_4_io_memIO_cen = iCache_io_SRAMIO_2_cen; // @[Top.scala 62:20]
  assign mem_4_io_memIO_wen = iCache_io_SRAMIO_2_wen; // @[Top.scala 62:20]
  assign mem_4_io_memIO_wdata = iCache_io_SRAMIO_2_wdata; // @[Top.scala 62:20]
  assign mem_4_io_memIO_addr = iCache_io_SRAMIO_2_addr; // @[Top.scala 62:20]
  assign mem_4_io_memIO_wmask = iCache_io_SRAMIO_2_wmask; // @[Top.scala 62:20]
  assign mem_5_clock = clock;
  assign mem_5_io_memIO_cen = dCache_io_SRAMIO_2_cen; // @[Top.scala 63:20]
  assign mem_5_io_memIO_wen = dCache_io_SRAMIO_2_wen; // @[Top.scala 63:20]
  assign mem_5_io_memIO_wdata = dCache_io_SRAMIO_2_wdata; // @[Top.scala 63:20]
  assign mem_5_io_memIO_addr = dCache_io_SRAMIO_2_addr; // @[Top.scala 63:20]
  assign mem_5_io_memIO_wmask = dCache_io_SRAMIO_2_wmask; // @[Top.scala 63:20]
  assign mem_6_clock = clock;
  assign mem_6_io_memIO_cen = iCache_io_SRAMIO_3_cen; // @[Top.scala 62:20]
  assign mem_6_io_memIO_wen = iCache_io_SRAMIO_3_wen; // @[Top.scala 62:20]
  assign mem_6_io_memIO_wdata = iCache_io_SRAMIO_3_wdata; // @[Top.scala 62:20]
  assign mem_6_io_memIO_addr = iCache_io_SRAMIO_3_addr; // @[Top.scala 62:20]
  assign mem_6_io_memIO_wmask = iCache_io_SRAMIO_3_wmask; // @[Top.scala 62:20]
  assign mem_7_clock = clock;
  assign mem_7_io_memIO_cen = dCache_io_SRAMIO_3_cen; // @[Top.scala 63:20]
  assign mem_7_io_memIO_wen = dCache_io_SRAMIO_3_wen; // @[Top.scala 63:20]
  assign mem_7_io_memIO_wdata = dCache_io_SRAMIO_3_wdata; // @[Top.scala 63:20]
  assign mem_7_io_memIO_addr = dCache_io_SRAMIO_3_addr; // @[Top.scala 63:20]
  assign mem_7_io_memIO_wmask = dCache_io_SRAMIO_3_wmask; // @[Top.scala 63:20]
endmodule
